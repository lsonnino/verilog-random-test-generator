`timescale 1ns / 1ps

`ifndef INSTR_MACROS
`define INSTR_MACROS 1

`define NO_INSTR 2'b00
`define WRITE_INSTR 2'b01
`define READ_INSTR 2'b10
`define MOVE_INSTR 2'b11
`endif

module testbench #(parameter DATA_WIDTH = 32, parameter BYTE_ADDR_WIDTH = 8, parameter BANKS_ADDR_WIDTH = 2);
    reg clk;
    reg rst;
    reg [1:0] op;
    reg [BYTE_ADDR_WIDTH+BANKS_ADDR_WIDTH-1:0] addr;
    reg [DATA_WIDTH-1:0] din;
    wire [DATA_WIDTH-1:0] dout;

    inspec uut (
        .clk(clk),
        .rst(rst),
        .op(op),
        .addr(addr),
        .din(din),
        .dout(dout)
    );

    initial begin
        $dumpfile("waveform.vcd");
        // $dumpvars(0, testbench.uut.rst, testbench.uut.op, testbench.uut.addr, testbench.uut.din, testbench.uut.dout);
        $dumpvars(0, uut);

        // Initialize
        clk = 0;
        rst = 1;
        op = `NO_INSTR;
        @(posedge clk); rst <= 0;
        @(posedge clk);

        // Autogenerated code        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h0, 8'h8a}; din <= 32'hfd33aafe;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h1, 8'h8a}; din <= 32'hf7a73d0e;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h2, 8'h8a}; din <= 32'hc57696f1;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h3, 8'h8a}; din <= 32'h7637746c;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h0, 8'h5e}; din <= 32'h18d88b97;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h1, 8'h5e}; din <= 32'h99b09031;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h2, 8'h5e}; din <= 32'h17e3a6ff;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h3, 8'h5e}; din <= 32'h954583ac;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h0, 8'h0b}; din <= 32'hb017d050;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h1, 8'h0b}; din <= 32'h28cd65bf;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h2, 8'h0b}; din <= 32'h33cfecea;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h3, 8'h0b}; din <= 32'hb97def85;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h0, 8'haf}; din <= 32'h2479e8b1;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h1, 8'haf}; din <= 32'hcdcc364c;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h2, 8'haf}; din <= 32'hfc7a10af;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h3, 8'haf}; din <= 32'hd150bc99;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h0, 8'h48}; din <= 32'heb892cda;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h1, 8'h48}; din <= 32'he52ecb82;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h2, 8'h48}; din <= 32'hf5eaace8;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h3, 8'h48}; din <= 32'hc3d97a77;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h0, 8'he4}; din <= 32'ha2f0179b;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h1, 8'he4}; din <= 32'h74feddfb;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h2, 8'he4}; din <= 32'h3ffb1d22;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h3, 8'he4}; din <= 32'h0c26ab5a;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h0, 8'h2d}; din <= 32'hbd29018b;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h1, 8'h2d}; din <= 32'h0b30f4aa;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h2, 8'h2d}; din <= 32'h53caf1d8;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h3, 8'h2d}; din <= 32'h2284bfe2;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h0, 8'h26}; din <= 32'h1a31d9ff;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h1, 8'h26}; din <= 32'h1bf93519;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h2, 8'h26}; din <= 32'h2ee0ac94;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h3, 8'h26}; din <= 32'h55d14d5a;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h0, 8'h50}; din <= 32'h58bbeb3f;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h1, 8'h50}; din <= 32'hf125f235;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h2, 8'h50}; din <= 32'h4740faa1;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h3, 8'h50}; din <= 32'h3f051834;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h0, 8'hc1}; din <= 32'h5a43d5cd;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h1, 8'hc1}; din <= 32'h6ebde513;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h2, 8'hc1}; din <= 32'h99904f8b;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h3, 8'hc1}; din <= 32'h814716b1;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h0, 8'ha6}; din <= 32'h0fb36ad3;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h1, 8'ha6}; din <= 32'h52e4da52;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h2, 8'ha6}; din <= 32'h3d4f96ce;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h3, 8'ha6}; din <= 32'h9ad56ea4;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h0, 8'he4}; din <= 32'ha4e1faf3;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h1, 8'he4}; din <= 32'h2c2208f4;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h2, 8'he4}; din <= 32'ha60c62a6;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h3, 8'he4}; din <= 32'hfdfb1767;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h0, 8'h87}; din <= 32'h37a110f6;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h1, 8'h87}; din <= 32'h37075aab;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h2, 8'h87}; din <= 32'h94810f51;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h3, 8'h87}; din <= 32'h4e4996f1;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h0, 8'h7c}; din <= 32'h1d80a715;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h1, 8'h7c}; din <= 32'hf1e64b9f;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h2, 8'h7c}; din <= 32'hb45b3719;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h3, 8'h7c}; din <= 32'hd7fc4091;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h0, 8'ha1}; din <= 32'he8340f6a;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h1, 8'ha1}; din <= 32'h1f57ffc5;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h2, 8'ha1}; din <= 32'h5b6f2754;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h3, 8'ha1}; din <= 32'h4fedd6af;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h0, 8'h00}; din <= 32'h696e0a41;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h1, 8'h00}; din <= 32'hafaadca8;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h2, 8'h00}; din <= 32'h4bf411a7;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h3, 8'h00}; din <= 32'h00d53ac5;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h0, 8'h6f}; din <= 32'hcdcddf58;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h1, 8'h6f}; din <= 32'hde50f92b;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h2, 8'h6f}; din <= 32'h2e6e32ff;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h3, 8'h6f}; din <= 32'h275dd17d;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h0, 8'he4}; din <= 32'h66151a22;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h1, 8'he4}; din <= 32'h8cc85f62;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h2, 8'he4}; din <= 32'hccac4211;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h3, 8'he4}; din <= 32'h4db66fb4;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h0, 8'h0b}; din <= 32'hc4474a9d;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h1, 8'h0b}; din <= 32'h553101e0;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h2, 8'h0b}; din <= 32'h58c2d28e;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h3, 8'h0b}; din <= 32'h1c1e30eb;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h0, 8'h94}; din <= 32'h01195662;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h1, 8'h94}; din <= 32'hd02efd69;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h2, 8'h94}; din <= 32'h25282091;
        @(posedge clk); op <= `WRITE_INSTR; addr <= {2'h3, 8'h94}; din <= 32'h74db2a69;

        // Finish
        @(posedge clk); op <= `NO_INSTR; addr <= 10'hxxx; din <= 32'hxxxxxxxx;
        repeat (5) @(posedge clk);
        $finish();
    end

    always #1 clk = ~clk;
endmodule
