`timescale 1ns / 1ps

module testbench #(parameter DATA_WIDTH = 32, parameter BYTE_ADDR_WIDTH = 8, parameter BANKS_ADDR_WIDTH = 2);
    reg clk;
    reg en, wen;
    reg [BYTE_ADDR_WIDTH+BANKS_ADDR_WIDTH-1:0] addr;
    reg [DATA_WIDTH-1:0] din;
    wire [DATA_WIDTH-1:0] dout;

    bank uut (
        .clk(clk),
        .en(en),
        .wen(wen),
        .addr(addr),
        .din(din),
        .dout(dout)
    );

    initial begin
        $dumpfile("waveform.vcd");
        // $dumpvars(0, testbench.uut.en, testbench.uut.wen, testbench.uut.addr, testbench.uut.din, testbench.uut.dout);
        $dumpvars(0, uut);

        // Initialize
        clk = 0;
        en = 0;
        wen = 0;
        @(posedge clk); en <= 0;
        @(posedge clk);

        // Autogenerated code        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c5; din <= 32'h504541e1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c7; din <= 32'hb43cc86f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h364; din <= 32'hfaa5d4b8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h097; din <= 32'hc601e54c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h206; din <= 32'h7363db64;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01c; din <= 32'h1602a02b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bc; din <= 32'h91f79e2b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h060; din <= 32'h29361a15;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15b; din <= 32'h819100b5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bc; din <= 32'heca1a885;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f0; din <= 32'h062407b0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h035; din <= 32'h8204f099;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0dd; din <= 32'h585f634c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04f; din <= 32'heab6a540;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04e; din <= 32'h3a18b770;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h006; din <= 32'h11dec3aa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d1; din <= 32'h201a3c2c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h009; din <= 32'h10d1041c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h338; din <= 32'h9eac28fe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f1; din <= 32'h2302b579;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h312; din <= 32'h11e24188;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h119; din <= 32'h03cd55b2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c2; din <= 32'h278f2977;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bb; din <= 32'hb368615f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31f; din <= 32'hc8d6f851;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h312; din <= 32'h388fb9f7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h392; din <= 32'h2df1d8de;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b1; din <= 32'ha221a4b5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20f; din <= 32'h24aa629c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h013; din <= 32'hdf2c909a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bb; din <= 32'haf51464d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h085; din <= 32'h976cc2f6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0eb; din <= 32'hb3b0152b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h334; din <= 32'hdeda348a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12e; din <= 32'h1d0d6a65;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c9; din <= 32'h2664758c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h337; din <= 32'h03cdce70;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11d; din <= 32'he33bc913;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d3; din <= 32'h9a133c85;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h330; din <= 32'hae54dbaa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h172; din <= 32'h6a8513e1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38c; din <= 32'hb2359350;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3dd; din <= 32'hbe99eac7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e1; din <= 32'h75f47204;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03a; din <= 32'hc0e58f50;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a0; din <= 32'h7ef223a9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h231; din <= 32'h8f56b911;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08a; din <= 32'he886d210;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h208; din <= 32'hdb0898fc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d5; din <= 32'h135e9f4a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26e; din <= 32'h17b1d787;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c4; din <= 32'he70e022c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h304; din <= 32'h4f494aaa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f1; din <= 32'h4342cdf7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h153; din <= 32'hff1a556a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a5; din <= 32'had315643;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ca; din <= 32'h6ead2b0d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27b; din <= 32'h0eccdda8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ac; din <= 32'h7f53447a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10b; din <= 32'h4a7ed39d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33c; din <= 32'h282edca7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h086; din <= 32'he528c22b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18a; din <= 32'h289fba2c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h019; din <= 32'hb8047295;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h089; din <= 32'h8fc6eb9f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ff; din <= 32'hf10ca0ed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15c; din <= 32'hda0c77a5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14e; din <= 32'hb53a404a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h181; din <= 32'h8c031c0b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h377; din <= 32'h3c46a41c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cb; din <= 32'he742acbc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22f; din <= 32'h1ffde76e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c1; din <= 32'h8e3208ee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h151; din <= 32'h0594387d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ab; din <= 32'h6384d841;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h237; din <= 32'h7ec49a50;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d7; din <= 32'h002811b6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h377; din <= 32'h258a652d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h265; din <= 32'hb45f1b60;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27f; din <= 32'hfd42dda7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ac; din <= 32'hf309746b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h234; din <= 32'h02eb129f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h253; din <= 32'h2f8ca253;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25e; din <= 32'h3dbb4b0a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h398; din <= 32'h75d7a043;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h025; din <= 32'h5e9c26e4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h346; din <= 32'h631cc722;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22b; din <= 32'h80e3b268;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d0; din <= 32'h1a1ccf6b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1df; din <= 32'h35b5131d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h083; din <= 32'hfc160f73;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h002; din <= 32'ha8892884;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h383; din <= 32'hbf991364;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e3; din <= 32'h3563bf61;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h288; din <= 32'h937aae60;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39f; din <= 32'h308655d2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34d; din <= 32'h4e9e5ecb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28e; din <= 32'ha7112462;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d2; din <= 32'h6229e62b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h388; din <= 32'hc9a83e3f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09d; din <= 32'hee506aed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h084; din <= 32'h53a906a7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h198; din <= 32'h1b896358;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h309; din <= 32'h4818b898;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24a; din <= 32'hcb912b3d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h345; din <= 32'h5c38c6d2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34b; din <= 32'h636ecc3b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h064; din <= 32'h133ce6c3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a7; din <= 32'h2bb3000a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39b; din <= 32'hb5f91af6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24a; din <= 32'h9601b663;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h260; din <= 32'hbecbffbe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fd; din <= 32'he24cc502;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3be; din <= 32'h8eeac3a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ff; din <= 32'h504e55b5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a5; din <= 32'h231f296d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fd; din <= 32'h3e41b803;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cc; din <= 32'h6605b0e9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fa; din <= 32'hdc02fba9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h190; din <= 32'he2d6fbe9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h273; din <= 32'he9995963;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d8; din <= 32'h492a44c3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h294; din <= 32'hb7dc5b57;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23c; din <= 32'h4fdcbe12;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h209; din <= 32'hf077584f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ba; din <= 32'h387724d5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h368; din <= 32'h09d538f7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d6; din <= 32'h0e880cf8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d4; din <= 32'h6bb22255;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d4; din <= 32'hb307a291;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h031; din <= 32'h05cae83d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33a; din <= 32'h7c610dbd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12a; din <= 32'ha80519f4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20f; din <= 32'h430fc78c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ae; din <= 32'h444a42ed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h262; din <= 32'hf6b5b910;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h281; din <= 32'hd0315c3d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h018; din <= 32'h149276b1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a9; din <= 32'hb60955b9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39a; din <= 32'h9ce0e911;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h322; din <= 32'h58f7e64a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cf; din <= 32'h94619aa9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e6; din <= 32'h4ec58dc3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2fe; din <= 32'ha2a4563b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h055; din <= 32'h24a95d9a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13c; din <= 32'h4c27a776;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a4; din <= 32'h403cd0f2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08a; din <= 32'hc467a712;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d4; din <= 32'h521422e5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h029; din <= 32'hc971a18e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bc; din <= 32'h374ff812;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a4; din <= 32'hb42a05a7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h287; din <= 32'h4d3bef88;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h349; din <= 32'h2158c6ff;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d7; din <= 32'h96edaf66;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h192; din <= 32'hc1c8a905;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h348; din <= 32'h88e6e2cc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f3; din <= 32'hab67c3ef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h029; din <= 32'haa1e58a1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05a; din <= 32'h17487e26;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ba; din <= 32'hafe2e5f5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h138; din <= 32'h2537932a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h315; din <= 32'h82ae3a07;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h005; din <= 32'hd4a8094f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e4; din <= 32'h33783be4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h088; din <= 32'h9c3ba5ca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h314; din <= 32'ha102f7c3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e4; din <= 32'h2574d445;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f9; din <= 32'hcf9ff2a5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26d; din <= 32'h6200550f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h257; din <= 32'hcd5c977a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cc; din <= 32'h740970ef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h277; din <= 32'hdc1f37b1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ac; din <= 32'h2f811c58;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a6; din <= 32'ha140d83b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h250; din <= 32'h4e03b6b6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2fe; din <= 32'ha3a90b4a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ce; din <= 32'hf4e60c69;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h058; din <= 32'h58e7132f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a7; din <= 32'h1c31cd62;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cb; din <= 32'h8d130a0d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33f; din <= 32'hc22239d8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h142; din <= 32'hddf208f2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37b; din <= 32'he09739ca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h236; din <= 32'h84afd735;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a2; din <= 32'ha462cd6a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h387; din <= 32'h9046934e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h284; din <= 32'h12d5f692;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bb; din <= 32'hbadf8838;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h196; din <= 32'he990c8f8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13b; din <= 32'h1748fdfa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h267; din <= 32'ha9a54ca9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h282; din <= 32'ha876190f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h076; din <= 32'hea23db0c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ef; din <= 32'hac4c412d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fb; din <= 32'hd571c70f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37a; din <= 32'h85372012;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ab; din <= 32'hbee274a4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11b; din <= 32'h0e2daecc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b2; din <= 32'h18a851ac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d5; din <= 32'h1c7e6361;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e7; din <= 32'h1e0767e5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h250; din <= 32'hc92ad4fe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d3; din <= 32'ha6372b24;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a2; din <= 32'h4e6a0800;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a9; din <= 32'he60610e3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1eb; din <= 32'h9c34c49c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e5; din <= 32'hf594e1a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h341; din <= 32'h161688f5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h164; din <= 32'hdccd7032;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h091; din <= 32'h9a8624f2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f8; din <= 32'h79f18544;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c8; din <= 32'hf00c9892;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h073; din <= 32'hcb7c27b9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39b; din <= 32'h983eb0b2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h263; din <= 32'h2895a4dc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10a; din <= 32'h3258fd58;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08c; din <= 32'h87edcc0d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h004; din <= 32'h23926ca7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h068; din <= 32'h7b9393c8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b8; din <= 32'h3769cb9d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38e; din <= 32'hadb87046;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26e; din <= 32'hd2723464;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10b; din <= 32'hb8bdde53;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13b; din <= 32'h3d5d6076;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e6; din <= 32'he1457aa5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h121; din <= 32'h80f21811;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h146; din <= 32'hb21e5c08;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h288; din <= 32'h1ccb868e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39d; din <= 32'h0d144507;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a7; din <= 32'h6886658b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37d; din <= 32'h04a178aa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bb; din <= 32'h8c65eca0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2da; din <= 32'h6f90a81d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05a; din <= 32'hfb4011b4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d2; din <= 32'h2056eaea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16e; din <= 32'hbda7b5d4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15e; din <= 32'hde65d9c5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33f; din <= 32'ha064b23d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12b; din <= 32'h07715413;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h082; din <= 32'h75f6f02a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1dd; din <= 32'h2fe2d61c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24d; din <= 32'h0e9d4a51;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h195; din <= 32'he52095a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h296; din <= 32'h09cfc709;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h248; din <= 32'he1c80b3d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h322; din <= 32'h0385a9f5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b6; din <= 32'h8251e30a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01c; din <= 32'hf83022fd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07d; din <= 32'hb525ee1e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h353; din <= 32'h813a0d83;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h317; din <= 32'he72f36dd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04d; din <= 32'h94eaadf6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c8; din <= 32'h97772abb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f5; din <= 32'hd31d42b7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h256; din <= 32'h7a53f7df;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b3; din <= 32'ha494992f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f5; din <= 32'h0633e061;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d4; din <= 32'hd054304b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h076; din <= 32'h2473a841;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a0; din <= 32'h71338841;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19f; din <= 32'h48031bfa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34e; din <= 32'h34f8e29e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h311; din <= 32'h38aec5c0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fa; din <= 32'hf4e2aab1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19c; din <= 32'hf331281d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h104; din <= 32'h9657c93b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e8; din <= 32'h829bf145;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h071; din <= 32'h5865cb9b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ea; din <= 32'h1d047c1c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h039; din <= 32'hf32a4195;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h057; din <= 32'he00024b8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h027; din <= 32'h87fb1a5b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h212; din <= 32'hb64b302f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08c; din <= 32'h8de4197b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h370; din <= 32'hed2e672d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d7; din <= 32'hc79dc579;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e1; din <= 32'hbc772400;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c5; din <= 32'h31c856ee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h188; din <= 32'h7dd5917c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f8; din <= 32'h2f89f25a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d1; din <= 32'h42028010;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ae; din <= 32'h33271d2f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h311; din <= 32'hc86e3da6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d7; din <= 32'h74914933;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h356; din <= 32'h7ff10e7b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h014; din <= 32'h39aeca93;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3dd; din <= 32'h2d15de2e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03e; din <= 32'h1757a592;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h103; din <= 32'hbc5dbc67;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h291; din <= 32'h5003286d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e7; din <= 32'h74d1a9c4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07b; din <= 32'h2de2e919;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23f; din <= 32'he83a2331;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c0; din <= 32'h3614a269;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d9; din <= 32'h3d2cebd1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f0; din <= 32'h80abb2cf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h073; din <= 32'h2dbf0eb9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h312; din <= 32'hc9c3b708;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21e; din <= 32'h15b83fac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e9; din <= 32'h06cfffc9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h153; din <= 32'hfbfe2dd4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17a; din <= 32'hab1e1ac4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d7; din <= 32'h2cf1c62a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36b; din <= 32'hfc56dcd8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03c; din <= 32'hb82d969e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h252; din <= 32'h4dfc2c4c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37d; din <= 32'hcbf0a8f7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ca; din <= 32'hdfbd97e1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h089; din <= 32'h0faa4368;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b9; din <= 32'h573ab810;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h144; din <= 32'h7f2d61c4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c2; din <= 32'h49948706;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18e; din <= 32'h893c5c39;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h191; din <= 32'h762ec74c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10a; din <= 32'ha68f39f0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h164; din <= 32'h5afb3a91;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16c; din <= 32'h436160fa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24d; din <= 32'hb1e48335;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h069; din <= 32'hf9457806;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h108; din <= 32'h7e50b290;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a2; din <= 32'head2d6e3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h353; din <= 32'h001ac915;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h275; din <= 32'h0b8a8080;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h217; din <= 32'h3b2d3cc9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h188; din <= 32'hb783f4a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h197; din <= 32'h5b7ae607;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h300; din <= 32'h60e90860;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a5; din <= 32'h6a819a21;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f4; din <= 32'h627f3f7a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e8; din <= 32'h332074d3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h206; din <= 32'h37dab9f0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h394; din <= 32'h3d9dde8e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h389; din <= 32'hfae594e9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ab; din <= 32'h2d01f3b6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26e; din <= 32'ha23100fa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e1; din <= 32'h90ba4761;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22c; din <= 32'hc02599a8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ce; din <= 32'ha759e9b9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a2; din <= 32'h4325a168;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h337; din <= 32'hfc97d923;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b1; din <= 32'h98d431c8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h378; din <= 32'h64303fa1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h325; din <= 32'hf41fa245;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h333; din <= 32'hd7a24f28;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h066; din <= 32'h0b8a531f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a3; din <= 32'h8d50b171;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h205; din <= 32'h3c5e2c7c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c2; din <= 32'h9f011053;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37d; din <= 32'h7dcbcdff;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h223; din <= 32'hd021c74b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e3; din <= 32'h98122010;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h019; din <= 32'h1cff0cfa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d9; din <= 32'hfeace1ad;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34f; din <= 32'h7685c473;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h261; din <= 32'h00639428;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f7; din <= 32'h106e2981;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h246; din <= 32'h9dd370f6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d3; din <= 32'h83b6eb50;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2db; din <= 32'hb6ba2859;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h265; din <= 32'h90a7e3d3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24f; din <= 32'ha1217314;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h093; din <= 32'h590ae527;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12b; din <= 32'h66c708b9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h174; din <= 32'ha32a3e37;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2aa; din <= 32'h595b69f0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33d; din <= 32'h68f66da7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h399; din <= 32'hfd7c02e0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h043; din <= 32'h4bdf476d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h220; din <= 32'h5e1b81b4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ab; din <= 32'h868618a5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bd; din <= 32'hb86f9708;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28f; din <= 32'hd170544e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e4; din <= 32'h08cfdcd3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h301; din <= 32'h2406949d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b0; din <= 32'h9c7947dd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14b; din <= 32'h9799cfd2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e4; din <= 32'hf140ff54;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h338; din <= 32'h61d64fd8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h170; din <= 32'hbc00b328;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h240; din <= 32'hf7b18b89;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b8; din <= 32'h63d0696b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04f; din <= 32'h3ca5fcda;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h060; din <= 32'hd2c4911f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h177; din <= 32'h4e2df988;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h093; din <= 32'hd6b70085;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ae; din <= 32'ha8ee0e3d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26f; din <= 32'h13465daf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h089; din <= 32'ha1e8bf2e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30a; din <= 32'h5aa47a87;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h132; din <= 32'h8900b1e5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d1; din <= 32'hfdf9bd85;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h116; din <= 32'hf3cbea59;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cb; din <= 32'h036c3d04;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h190; din <= 32'h247611cb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2eb; din <= 32'hb3294556;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h204; din <= 32'hd5949133;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1de; din <= 32'h33ea4b4c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e5; din <= 32'h05933c0e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h127; din <= 32'h113e912d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h130; din <= 32'hda4a9b8d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09d; din <= 32'h8b08cc3e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ea; din <= 32'h5c51f3be;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d0; din <= 32'hdc870d52;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h335; din <= 32'had32a4ad;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h376; din <= 32'h1c0b4549;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h176; din <= 32'h52c4241a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h055; din <= 32'h9def8f43;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f2; din <= 32'h97d2b6af;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cb; din <= 32'h50df34c3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21c; din <= 32'ha15d846a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h272; din <= 32'he823f928;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h209; din <= 32'h45948fea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06d; din <= 32'hb6439eb2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h253; din <= 32'h99decd8a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h045; din <= 32'h3416497a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h075; din <= 32'h327ada75;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06a; din <= 32'h13a00fa3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h345; din <= 32'h5a1524ce;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h068; din <= 32'h12edb41f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27f; din <= 32'hde123158;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15d; din <= 32'h64524913;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17f; din <= 32'hc51d3eb0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d5; din <= 32'ha94c4dcd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cb; din <= 32'h6ea57481;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fb; din <= 32'hde0a7a20;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c5; din <= 32'hda7c62c0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h232; din <= 32'hf070c710;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h252; din <= 32'h02a732bd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2fe; din <= 32'hebf5176c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h088; din <= 32'h137af9ca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b3; din <= 32'hf886f5f3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a7; din <= 32'h8056c47a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h398; din <= 32'h678f563c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b5; din <= 32'hcf26b110;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36f; din <= 32'hf97ddb22;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19e; din <= 32'hdc2dc16a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h237; din <= 32'hea5839cc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c8; din <= 32'hae989d01;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b8; din <= 32'h3d401c34;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h160; din <= 32'h98485591;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h383; din <= 32'h5d561edd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b9; din <= 32'h328cb2cb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ee; din <= 32'ha0144940;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ec; din <= 32'ha2766070;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17e; din <= 32'hacb45043;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16e; din <= 32'h43a8c7eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h170; din <= 32'h220a8ba2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h181; din <= 32'h6904a764;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bd; din <= 32'hfbc5050d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h236; din <= 32'h2ce29bba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26f; din <= 32'ha42c7946;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06d; din <= 32'h9bda82db;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f2; din <= 32'hac5d8efd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h053; din <= 32'h0a940404;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h034; din <= 32'hd14b6281;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h134; din <= 32'hea92bb0b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28c; din <= 32'h38e32519;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24c; din <= 32'h1102aac6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f8; din <= 32'hba799d45;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h356; din <= 32'h98e77b4d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h017; din <= 32'h3d5dc789;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25b; din <= 32'h615ae69a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ac; din <= 32'h88ea16c6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h359; din <= 32'hb6afbd17;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ed; din <= 32'hf27c80ce;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h283; din <= 32'h501efb4f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a7; din <= 32'h6317ee84;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e6; din <= 32'h5cea9c81;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h147; din <= 32'h942e0c30;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2fe; din <= 32'h8b6683a7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h136; din <= 32'h2f2fe713;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h281; din <= 32'h10f10474;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e5; din <= 32'h92dca5ee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h039; din <= 32'h2e794394;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h040; din <= 32'hff6b4adb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h066; din <= 32'h898b167e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24b; din <= 32'h0871cf1e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35d; din <= 32'ha92a5e34;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h246; din <= 32'hc64c30c2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h037; din <= 32'h55e74dc0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h104; din <= 32'h433f6e8a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h134; din <= 32'h517335d7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bc; din <= 32'h5345bfb2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cc; din <= 32'h8fe58124;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h134; din <= 32'hfb81d583;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h250; din <= 32'h3889b293;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ef; din <= 32'h12b372ea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c4; din <= 32'h60e6141a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h174; din <= 32'h3d480a19;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h122; din <= 32'h6f749803;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14e; din <= 32'h642fab23;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h249; din <= 32'hd221a2fb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b6; din <= 32'h379d1638;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c1; din <= 32'he833092d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h294; din <= 32'hc0cae475;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22c; din <= 32'h1048065a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15e; din <= 32'hd28127c3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h396; din <= 32'hd48f1511;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c3; din <= 32'he92fc9a2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c8; din <= 32'hd25afa30;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08c; din <= 32'hd42ef17c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h227; din <= 32'h4d037427;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h060; din <= 32'hcc4c158b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h220; din <= 32'hffc24b3e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23d; din <= 32'hf3d296ac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e3; din <= 32'h6d7de64f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h049; din <= 32'hb9b2798d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h039; din <= 32'h7abd03db;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h094; din <= 32'h55dc7e3b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h173; din <= 32'h7013d282;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h346; din <= 32'hedf46be5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h328; din <= 32'ha77adf19;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a6; din <= 32'h67abfa5e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h341; din <= 32'ha0ad18c7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20e; din <= 32'h1ef76989;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e1; din <= 32'hb10c2c53;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bf; din <= 32'h9eac91e2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e3; din <= 32'h91081c18;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e3; din <= 32'h658c91b8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27d; din <= 32'h01cf2f11;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h349; din <= 32'h33cf698d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h169; din <= 32'h55d476ab;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c0; din <= 32'h620411e8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08f; din <= 32'h0f887c82;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1de; din <= 32'h158b409f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36f; din <= 32'h78b56e55;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h390; din <= 32'hda7f761e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fe; din <= 32'h398150e7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h285; din <= 32'h4145dade;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1da; din <= 32'h980a0e21;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h279; din <= 32'hb7120b33;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h241; din <= 32'hf850bda0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35f; din <= 32'h8a26cda6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19d; din <= 32'h9cfcb1b3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08b; din <= 32'hc166b949;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f1; din <= 32'hf691f876;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25c; din <= 32'h62effd99;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h265; din <= 32'he7619d9c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h051; din <= 32'ha54b6db7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h155; din <= 32'h9d72cc4e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15e; din <= 32'hc6cf21ad;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3de; din <= 32'h94ed77db;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f2; din <= 32'h237005e3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c5; din <= 32'h870ec14e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h249; din <= 32'h009a64d7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h005; din <= 32'h2a1ae8cc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13c; din <= 32'h969b08f5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h125; din <= 32'hd1a26ea0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h090; din <= 32'ha63a7eb4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e1; din <= 32'hc1a29bc3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h070; din <= 32'ha70540ba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h078; din <= 32'h6da746c8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11f; din <= 32'h1c9b8046;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h185; din <= 32'he821b63e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h381; din <= 32'hf4bfa2b5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h392; din <= 32'h6307a7d7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fd; din <= 32'h5663fa19;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ba; din <= 32'h1e4707e6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h292; din <= 32'h27eab25f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fb; din <= 32'he6953f71;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b5; din <= 32'hef2bbec8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h289; din <= 32'hb07c4100;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e4; din <= 32'hb97fa496;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05d; din <= 32'h4b2a0d0b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h205; din <= 32'hd1c7a83b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h388; din <= 32'h8477bb58;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h045; din <= 32'h7386de2a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h233; din <= 32'h2ecdfa41;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h240; din <= 32'hd5fe5c78;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2dc; din <= 32'haa2e1f45;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h252; din <= 32'hee55939b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d6; din <= 32'heeda6761;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a3; din <= 32'h2a75e728;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11c; din <= 32'h5a8aaee6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h050; din <= 32'h44829c45;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a2; din <= 32'h68739257;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11d; din <= 32'hd99b4fa9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ae; din <= 32'h0c1852e1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d5; din <= 32'h5d870d51;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a6; din <= 32'h97e1dbb2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h146; din <= 32'h479ee2a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05e; din <= 32'h17274a08;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0dc; din <= 32'h634941c9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h283; din <= 32'h77d8681e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26b; din <= 32'ha1a239ce;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c3; din <= 32'he0645575;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21a; din <= 32'hb48f9aed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h287; din <= 32'h6dde5616;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h048; din <= 32'hefe5904a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h359; din <= 32'h8a0cded4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05d; din <= 32'hb8904c91;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a2; din <= 32'h0af6ba41;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h371; din <= 32'hcdabe3ca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d0; din <= 32'ha7098c3f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1dd; din <= 32'h535d9ef4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h157; din <= 32'h315a7b21;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h157; din <= 32'h57efb006;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a4; din <= 32'h3c7171c5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ec; din <= 32'hf5702585;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22e; din <= 32'h5e5bcc9e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a6; din <= 32'head9530a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h055; din <= 32'h2ed0e85d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37c; din <= 32'h342f9c0f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cf; din <= 32'hf937a1db;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h294; din <= 32'he12390df;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22a; din <= 32'habc9c844;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3af; din <= 32'h3ae70684;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h050; din <= 32'hf7a178af;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h015; din <= 32'hb2e84cae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h391; din <= 32'h72357ac5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d4; din <= 32'h02a74981;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h083; din <= 32'h6388ccdc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h391; din <= 32'h4904698c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a9; din <= 32'h7c42a67c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20a; din <= 32'h7d539dae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24f; din <= 32'h0dc8291b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0af; din <= 32'ha658fb3a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09d; din <= 32'ha9a7090d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ac; din <= 32'hac402a9d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31f; din <= 32'h59bf3654;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35f; din <= 32'h61202970;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28a; din <= 32'h0d5f87cf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b2; din <= 32'h9ad835cd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h191; din <= 32'h09b8ebf0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04d; din <= 32'h28232cf8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13e; din <= 32'ha2a2fcc9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2be; din <= 32'h0b81ead6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f4; din <= 32'h79c88bdc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38a; din <= 32'hc61102a9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01e; din <= 32'h86ca3f7f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31f; din <= 32'hcfc82286;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h138; din <= 32'hfd9d5638;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27e; din <= 32'he009abd8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h250; din <= 32'h39dfe79a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17c; din <= 32'h5bc74e99;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h127; din <= 32'h0e9e541f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h085; din <= 32'h29aa8c59;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h268; din <= 32'hd042b7aa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ab; din <= 32'hbc9c7300;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h012; din <= 32'h1326c150;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h122; din <= 32'h90a444d5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a4; din <= 32'h7b63ae77;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h108; din <= 32'hd8e62762;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h173; din <= 32'hd5dd5a18;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06f; din <= 32'h18358fad;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h052; din <= 32'h23bc5595;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d1; din <= 32'hbae09386;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09f; din <= 32'heb529a33;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h347; din <= 32'h244170ef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08a; din <= 32'hba5b746a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e5; din <= 32'h68dabe30;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d9; din <= 32'h02df2f36;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h273; din <= 32'h42703ce9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h174; din <= 32'habe67a5a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32c; din <= 32'hcae6fec8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h273; din <= 32'he9e44fc8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h065; din <= 32'h70c4a1d2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h130; din <= 32'hd734fcc9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h161; din <= 32'h6fc9c105;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h320; din <= 32'h9e7ae5ca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h351; din <= 32'h6f1d98f5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24c; din <= 32'h07113fb1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cf; din <= 32'h57600c5d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e0; din <= 32'h540400b5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h234; din <= 32'h2601cc69;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h196; din <= 32'hcb5c24ac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39a; din <= 32'h034e43d2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09b; din <= 32'h6bb5974f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b8; din <= 32'hccb3daba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h008; din <= 32'hd20a241d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27d; din <= 32'hef11e67b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h029; din <= 32'ha062e800;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bb; din <= 32'h8b47f185;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ea; din <= 32'h7196e2f2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34f; din <= 32'hd0b8d6bd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h303; din <= 32'h96116ce4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h303; din <= 32'hce6983cf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0dc; din <= 32'ha080b015;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h070; din <= 32'heeada820;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38a; din <= 32'h03188e34;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f4; din <= 32'h39230354;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ad; din <= 32'hbb2a604a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h153; din <= 32'h832ba860;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h177; din <= 32'h5e7aaa3d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25a; din <= 32'h5bcdffaa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18c; din <= 32'hfc8ad489;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h317; din <= 32'hb02ab594;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h169; din <= 32'h7febeef2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h204; din <= 32'hd0de7ed4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h103; din <= 32'hd2a22182;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b4; din <= 32'ha2f729c7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c0; din <= 32'h3cfcffd2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h251; din <= 32'ha4a92c4a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b9; din <= 32'hf6b0388c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cd; din <= 32'h8f5f97ce;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h210; din <= 32'haf3c15d9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20a; din <= 32'h8d823f44;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30a; din <= 32'h114d5cff;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36c; din <= 32'hcba886b8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39a; din <= 32'hd12d0c6b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28d; din <= 32'h5e54864c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a2; din <= 32'h59e9c87a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h346; din <= 32'h6881f91b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f0; din <= 32'h2dfc70b2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a7; din <= 32'hf45d3bc1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14a; din <= 32'hca5641a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h009; din <= 32'h59affb8b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h054; din <= 32'h126c3b10;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d8; din <= 32'h0723f64d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h163; din <= 32'h295c2d89;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h194; din <= 32'he8e9554f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h274; din <= 32'h3eceab7e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04a; din <= 32'h111000c5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20f; din <= 32'h1cf6d34f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e9; din <= 32'hf9651d7a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h132; din <= 32'ha72a8aac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h125; din <= 32'h97d94013;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h125; din <= 32'hafb43a7c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h275; din <= 32'h06829422;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c8; din <= 32'h0becaef4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h251; din <= 32'h768ce8ab;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h112; din <= 32'h8b1e0b1e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h195; din <= 32'h0329852b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h111; din <= 32'h6af91e0a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d1; din <= 32'h806d26a8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21d; din <= 32'h64fc07ca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12b; din <= 32'ha29c029e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e6; din <= 32'h9c9986f9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38a; din <= 32'h5cdebb9a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h302; din <= 32'h4b5dc3f4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f8; din <= 32'h6d700843;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bb; din <= 32'hf5564297;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0dc; din <= 32'h22024dae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h049; din <= 32'h80f55d0a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a3; din <= 32'h4f60dd8c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a8; din <= 32'h8e866f12;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bc; din <= 32'h096409c6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e3; din <= 32'h6d7f96f6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cd; din <= 32'h5e6f0543;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h398; din <= 32'h63ac7faa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23c; din <= 32'hc06b1b0e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21f; din <= 32'hc932f299;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h256; din <= 32'h280a9d49;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h247; din <= 32'he7769994;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37f; din <= 32'hae16744f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a0; din <= 32'h5a56a520;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36e; din <= 32'h2de5cda4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h181; din <= 32'h31ed7073;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ad; din <= 32'h8d0988fb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d2; din <= 32'h3982f842;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25b; din <= 32'h5ff2a6f4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03e; din <= 32'h5b14a468;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bf; din <= 32'hb6d78f4f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h065; din <= 32'hac87a849;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26f; din <= 32'h5b724894;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bc; din <= 32'hc2bc0084;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e9; din <= 32'h9793de6f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34d; din <= 32'h5c576e20;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13a; din <= 32'hb988a486;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h251; din <= 32'h74c4fa36;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h038; din <= 32'hb25cc77b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2fc; din <= 32'h6d2cbd74;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06f; din <= 32'h3519c34f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31b; din <= 32'h093b41e5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f8; din <= 32'h64ff1468;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h075; din <= 32'he08521fb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17a; din <= 32'hfdba3924;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h000; din <= 32'h1b5a2ec2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e1; din <= 32'h641d1394;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08d; din <= 32'h7375a3f0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h206; din <= 32'h95dbb4ec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h100; din <= 32'he3d98b09;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e9; din <= 32'h8e17b643;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1db; din <= 32'h449da87e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h064; din <= 32'hcfc83e79;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d4; din <= 32'ha7461089;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h320; din <= 32'hadc934fd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25e; din <= 32'h3f8e7b0c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h304; din <= 32'hc595271b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37a; din <= 32'h95aa7db1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h014; din <= 32'hd206db28;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h351; din <= 32'h13498b8e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cf; din <= 32'hd4874cd4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h130; din <= 32'h913dc2a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b0; din <= 32'h213fc072;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bf; din <= 32'hfd6e358f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h169; din <= 32'h096eabb8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a7; din <= 32'h01d6ec17;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h036; din <= 32'h4de03c9c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ed; din <= 32'hd5bb0b28;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1aa; din <= 32'h07e14f90;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h000; din <= 32'h971ca1a5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16d; din <= 32'hac98f714;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fb; din <= 32'h6ed0d26e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f3; din <= 32'h8914795c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ff; din <= 32'h47cce6ed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b5; din <= 32'h54155b99;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h380; din <= 32'ha516c529;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h238; din <= 32'h16fd2d17;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f6; din <= 32'h435719d4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fb; din <= 32'h13f6925d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e5; din <= 32'h310b3d08;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h095; din <= 32'h5e93d719;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ce; din <= 32'h6d85ba4c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h379; din <= 32'hd6205309;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h266; din <= 32'he324fbfe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f2; din <= 32'h9e6235a4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h137; din <= 32'hd39961c8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08c; din <= 32'h9e356d12;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h343; din <= 32'hd2cf5902;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a8; din <= 32'hd0693c14;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e3; din <= 32'h1abd32fa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h070; din <= 32'hbb516484;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h165; din <= 32'hc8e6cf22;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c7; din <= 32'ha8f5195d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h101; din <= 32'he06cf259;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h216; din <= 32'h2ab083fc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h393; din <= 32'h0d5e5c2c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h145; din <= 32'hc7c4decf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10a; din <= 32'h9abc110d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h291; din <= 32'hdf1f7ebb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20c; din <= 32'h99e5d015;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c6; din <= 32'h3a088378;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h364; din <= 32'hcfec9312;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c7; din <= 32'hf6f5e1b1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f1; din <= 32'hff2e5af8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h153; din <= 32'he3fc8c65;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1de; din <= 32'h56ba6d60;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00f; din <= 32'h391ea8f4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26f; din <= 32'h5782e9cd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ee; din <= 32'h66fa920f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h353; din <= 32'hf5bfad65;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h059; din <= 32'h063b327d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h161; din <= 32'h8eda50ac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d3; din <= 32'h898b3559;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27a; din <= 32'h8b3b8fec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h048; din <= 32'hb384b75c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fc; din <= 32'h33883042;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h245; din <= 32'hf928edd3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h266; din <= 32'h69f10642;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h338; din <= 32'h2134accf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h393; din <= 32'h1a09d145;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33c; din <= 32'h75de9619;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h313; din <= 32'hd7498175;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07d; din <= 32'h193b0c4f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20e; din <= 32'h19482b5b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c1; din <= 32'h3cde6916;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22e; din <= 32'h84f65b85;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h148; din <= 32'h53ff5065;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h117; din <= 32'hb02d077e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h380; din <= 32'h8a4e26ff;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1de; din <= 32'h8624c541;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0be; din <= 32'haf33f422;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h044; din <= 32'hd935011e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h306; din <= 32'hf9a6c771;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f3; din <= 32'h8241fd1d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2db; din <= 32'h69bc79eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h093; din <= 32'hc0fdac66;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16c; din <= 32'h98f26569;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h154; din <= 32'h8de3ef9e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c1; din <= 32'h20adfd4d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h339; din <= 32'h7bd1a025;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17b; din <= 32'hb23bc418;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d6; din <= 32'h520ce925;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h251; din <= 32'h41f6dafd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fb; din <= 32'h38606b1a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f0; din <= 32'hc8faeb4e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h373; din <= 32'h015f7bae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a7; din <= 32'hb093af8a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07d; din <= 32'hab19a656;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c7; din <= 32'h349c5ede;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h154; din <= 32'h7851d08e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16d; din <= 32'h2e2fdc89;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h335; din <= 32'hd88ce6f3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26c; din <= 32'h7a16bbab;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h213; din <= 32'h6db2cc7d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ca; din <= 32'h6a848bc2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34b; din <= 32'hc1d7885d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cd; din <= 32'h00732bb7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f7; din <= 32'h3556ff8f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06f; din <= 32'h374313a5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25e; din <= 32'h8dbd6a20;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h051; din <= 32'hc2174af8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2fa; din <= 32'h447b6da8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20b; din <= 32'hbea8e647;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bf; din <= 32'hfac0dac1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f2; din <= 32'h5de4dabd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f6; din <= 32'h31ec536b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00c; din <= 32'h77e7113d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h189; din <= 32'h5800b74a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h120; din <= 32'hd1d371ae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e7; din <= 32'h559a47dd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h172; din <= 32'h9919bc59;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h345; din <= 32'hebdfc416;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c3; din <= 32'h241b6458;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b4; din <= 32'h585d9f00;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b5; din <= 32'h6a5c2bc1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e6; din <= 32'h8b03adf3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h364; din <= 32'h494b8ab8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02a; din <= 32'h5045dc1e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h115; din <= 32'h22fa0db5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ed; din <= 32'h597b0386;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25c; din <= 32'hcf9e45c7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2eb; din <= 32'h51f06810;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h205; din <= 32'hc8793dac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05b; din <= 32'h8bce5537;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h018; din <= 32'h058dbc21;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fd; din <= 32'ha288b5ec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fb; din <= 32'h1fa0a754;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h049; din <= 32'h10c52888;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bb; din <= 32'hd8cb588b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h089; din <= 32'h3740edb3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h316; din <= 32'hb2f3af5d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12d; din <= 32'hae2f90cb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3df; din <= 32'heee4555f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39e; din <= 32'h0e89778b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h340; din <= 32'h0338bd97;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h354; din <= 32'h097e6830;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17f; din <= 32'h4521c076;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c4; din <= 32'h269a0900;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h297; din <= 32'hc37cc069;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cc; din <= 32'hdfeac298;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05f; din <= 32'hd786efe7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0eb; din <= 32'ha10a8ffe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h150; din <= 32'h0cf03481;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ea; din <= 32'h27127014;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h110; din <= 32'hd4b90956;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h258; din <= 32'h8662a429;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c9; din <= 32'h87d04fe9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29c; din <= 32'hc5383ec1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h368; din <= 32'h9d34e822;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f2; din <= 32'h4725d974;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2db; din <= 32'h326f78f8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21a; din <= 32'h82e72180;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h025; din <= 32'h45097437;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09b; din <= 32'hdf3344a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b2; din <= 32'h06cf6fb6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h103; din <= 32'h78bda362;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ec; din <= 32'h0f7cb352;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h067; din <= 32'h16379df8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20d; din <= 32'h313fc4b6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h327; din <= 32'h0d53a5a5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37f; din <= 32'h399fd419;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h376; din <= 32'h2d124a60;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2eb; din <= 32'h372b1891;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a2; din <= 32'hbe8b10a7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h262; din <= 32'hc69a252d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d8; din <= 32'h25fc1afa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09a; din <= 32'h78cbcf1b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f3; din <= 32'h608e5989;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bf; din <= 32'h07763c8a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h073; din <= 32'hb43ef6cb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37b; din <= 32'h71d3de0f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a9; din <= 32'h79cf6dfc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h187; din <= 32'h52104b3c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1aa; din <= 32'h7c97c211;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03d; din <= 32'hfa7805a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13f; din <= 32'h6594cc34;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14b; din <= 32'h48a40400;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24d; din <= 32'h1908fba6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h178; din <= 32'hcff3d70b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04c; din <= 32'h03596e76;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h009; din <= 32'hb640c1b2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h254; din <= 32'h7a789cca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h017; din <= 32'h5ae39fa3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19d; din <= 32'hf204f89e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h189; din <= 32'h7b099f10;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1dd; din <= 32'he385da55;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ce; din <= 32'h3ca02d2a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00c; din <= 32'h78ef79c0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ea; din <= 32'hd11ebc32;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d1; din <= 32'hc59575a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a1; din <= 32'h72df5aa1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h086; din <= 32'hb242cba0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16e; din <= 32'heae7fe49;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h081; din <= 32'hb5bfff70;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a6; din <= 32'h6e228665;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b8; din <= 32'h945c3c0f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b7; din <= 32'h2f24c37f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ea; din <= 32'h68f9aa6e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h233; din <= 32'h8a934ed8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10a; din <= 32'h587231a1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02f; din <= 32'h7e4169c7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f6; din <= 32'h7e3d8052;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01f; din <= 32'hfad98364;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21a; din <= 32'h80f91f2e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c6; din <= 32'h86cc9f12;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h290; din <= 32'h42c8bf71;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f2; din <= 32'h15e46185;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13e; din <= 32'hc97e8c9b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bd; din <= 32'h2f083467;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35d; din <= 32'hb509a30a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h300; din <= 32'h0b097300;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1df; din <= 32'hdb968030;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c9; din <= 32'h73507aee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15d; din <= 32'h6a691a3c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h039; din <= 32'h45d80a16;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ac; din <= 32'h43b12b5e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h301; din <= 32'hac362648;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h076; din <= 32'he33e3608;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f8; din <= 32'ha91f7fd2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ba; din <= 32'h1790d072;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36f; din <= 32'h4c836178;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ca; din <= 32'hd3f48d21;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h233; din <= 32'h10daf669;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04e; din <= 32'h9e1b57d6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e8; din <= 32'h8fe9e1fa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b6; din <= 32'h4f17f1a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b6; din <= 32'h5af7b8f7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a5; din <= 32'h5ad24778;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f5; din <= 32'h35c4320c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a7; din <= 32'h6301b7d2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31c; din <= 32'h6c3a0881;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h079; din <= 32'hc7a0aa86;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a4; din <= 32'h384e2299;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h092; din <= 32'hd2f86cc8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h106; din <= 32'h44cfebaa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h387; din <= 32'h88d3edf4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37c; din <= 32'hed8f3726;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ac; din <= 32'he65a058a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bb; din <= 32'h4937925a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h278; din <= 32'hb2a850bf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09e; din <= 32'h680ed4a1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01b; din <= 32'ha56043b1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23b; din <= 32'h9f53628e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31b; din <= 32'h78c63e00;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b1; din <= 32'h7b24951c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h203; din <= 32'h5da0978c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ac; din <= 32'h3c3c9caf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e5; din <= 32'h60d9136a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11c; din <= 32'h45778624;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24a; din <= 32'h6d8c0f86;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f5; din <= 32'hea172fb8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h398; din <= 32'h3b9232eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h061; din <= 32'h685472c3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f6; din <= 32'hef4534f9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c8; din <= 32'h34243ab6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h329; din <= 32'h95ced0aa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c7; din <= 32'hbdf13c57;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f8; din <= 32'h3bbedcf0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h023; din <= 32'h033aa578;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b1; din <= 32'h1af1f469;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h284; din <= 32'he5fa1570;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h019; din <= 32'hceae9493;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h072; din <= 32'h8b13b037;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h180; din <= 32'hf744be15;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h359; din <= 32'h2ff294ca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e8; din <= 32'hd7042c84;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33d; din <= 32'h0e5ebcb3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h197; din <= 32'h91968fe6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h343; din <= 32'h390f6834;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b8; din <= 32'hd575e73b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h246; din <= 32'hfa2a9086;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ef; din <= 32'hf1721737;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31e; din <= 32'hbb4a2817;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a8; din <= 32'hb7b17824;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e1; din <= 32'h089e6133;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h396; din <= 32'h1ca93f48;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h051; din <= 32'h0f5c632e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h182; din <= 32'hf6aacdaa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a3; din <= 32'hcf6faea1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c4; din <= 32'he077a932;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h307; din <= 32'hf5db0386;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h078; din <= 32'h2d019043;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02b; din <= 32'h31024c49;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c8; din <= 32'h4ae656cc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h217; din <= 32'h7f0235a4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h338; din <= 32'h2ecad0a4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20d; din <= 32'h4071dde6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fe; din <= 32'ha5a78948;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bc; din <= 32'hcb6124f3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22e; din <= 32'h598efcdf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bc; din <= 32'hdfcf5f3f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30e; din <= 32'h19c2fa60;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h223; din <= 32'h4a4614da;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d7; din <= 32'habf32081;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c1; din <= 32'h1c7c6422;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c2; din <= 32'h6578aeeb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a4; din <= 32'hb84759a1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h038; din <= 32'h7a23ff91;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3dd; din <= 32'h452d18af;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32d; din <= 32'heea9cff5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21e; din <= 32'h661eebce;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38d; din <= 32'h6b906126;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h081; din <= 32'h81acb95d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h209; din <= 32'h088ebf70;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09e; din <= 32'hc5ddd43c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ca; din <= 32'h7b0f2b88;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ce; din <= 32'h6fbffaef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ca; din <= 32'h0e53e247;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h265; din <= 32'hdf5399ec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h174; din <= 32'h1939b995;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27c; din <= 32'h26a369b9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16c; din <= 32'hcf4e4e16;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h034; din <= 32'h98977e1c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23d; din <= 32'h1a4ab522;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a9; din <= 32'h3c494cb8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fc; din <= 32'h79705628;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b1; din <= 32'h320d803d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h351; din <= 32'hbb428e1e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h389; din <= 32'h4f0803ca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h156; din <= 32'h5092d6c8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3de; din <= 32'hae1e74f3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h271; din <= 32'h90b65e2a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25f; din <= 32'h8a10791b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d3; din <= 32'hc9225ebf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h212; din <= 32'h56d722eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23b; din <= 32'h4452e926;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33f; din <= 32'hb496b979;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39c; din <= 32'h63374c5e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34d; din <= 32'h2e364ee3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h378; din <= 32'h9d5240a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d5; din <= 32'h38e607d4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a0; din <= 32'ha018d311;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26e; din <= 32'h4399008b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c6; din <= 32'h5b2b73cf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0db; din <= 32'h73267fe7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h394; din <= 32'h957a30a7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36f; din <= 32'h7c6b775e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ad; din <= 32'h43c7133e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36e; din <= 32'hf73948b0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h068; din <= 32'h826ad61d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06e; din <= 32'h268a8b98;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f7; din <= 32'he9ce94b6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1eb; din <= 32'h95482476;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39c; din <= 32'hb37fbfb9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h055; din <= 32'h3c6df468;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h325; din <= 32'ha65a08a1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02a; din <= 32'h0a3f0455;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28e; din <= 32'h486b41ec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a7; din <= 32'hb035bec9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ee; din <= 32'hf1552732;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h002; din <= 32'h5fc8bdea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f0; din <= 32'h92499a95;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0db; din <= 32'h91b0b7b8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h214; din <= 32'hb52ddae6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d8; din <= 32'h690f9584;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ba; din <= 32'h4d420969;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04a; din <= 32'h84a27725;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38a; din <= 32'he7a7a817;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05a; din <= 32'hfc835cca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0eb; din <= 32'h5dadbe97;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a4; din <= 32'hbb1bb0b3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28c; din <= 32'ha1c88db1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d3; din <= 32'h2792437a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h172; din <= 32'he16aa524;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h189; din <= 32'h2fa413b8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14e; din <= 32'h58a0220e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15d; din <= 32'h3b7b19cd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b2; din <= 32'h4b377fff;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28b; din <= 32'h9906ea58;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h327; din <= 32'h39ff8c29;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3db; din <= 32'h918273ad;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d8; din <= 32'hd8ff8e08;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cf; din <= 32'ha7c77c84;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c2; din <= 32'h83dd23ba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h353; din <= 32'h5ce893f9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00e; din <= 32'hfc7a8eab;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ad; din <= 32'h3a15350c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19f; din <= 32'h28a33ede;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h144; din <= 32'hbdd1f61a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h298; din <= 32'h45604303;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d8; din <= 32'h66385cda;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36f; din <= 32'haedc5c95;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h345; din <= 32'h250cce91;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26c; din <= 32'ha60e94d9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e5; din <= 32'h73139547;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c7; din <= 32'h2702b4cc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h077; din <= 32'h580eea94;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h279; din <= 32'h52380080;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h225; din <= 32'h748faf8e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29b; din <= 32'hac9d9144;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cb; din <= 32'h02b6ec88;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bc; din <= 32'hd284b400;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h125; din <= 32'hc2a7e8a8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h397; din <= 32'hee7f5bc2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h082; din <= 32'h0c905505;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h022; din <= 32'h91b474f5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a9; din <= 32'hb4faec1a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h026; din <= 32'h5b9f6c05;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h179; din <= 32'h86ea44ad;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37d; din <= 32'h96e2e821;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h331; din <= 32'h5018bde0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2eb; din <= 32'hbe1c3a7f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h092; din <= 32'h4ba86fe7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28c; din <= 32'he5a5b104;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h034; din <= 32'h8a0f6642;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h363; din <= 32'h0a062516;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a6; din <= 32'h05713996;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24d; din <= 32'ha19601e3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d6; din <= 32'hf7185297;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bf; din <= 32'h03d8d5a2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ee; din <= 32'hf43c0ed5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cd; din <= 32'hf790a67d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17c; din <= 32'ha1fcd750;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h126; din <= 32'hbce4f589;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d3; din <= 32'hcffcd816;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c1; din <= 32'h83da8520;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a9; din <= 32'h976c4583;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20f; din <= 32'h27a09753;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d1; din <= 32'h40c12781;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h055; din <= 32'h508a01e6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a7; din <= 32'h5ab99419;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36e; din <= 32'h8045c805;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h201; din <= 32'h4a31b593;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e7; din <= 32'hc7257fc4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36f; din <= 32'h9060cd9c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27c; din <= 32'h9ad70847;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h213; din <= 32'hfdb7ab6b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24d; din <= 32'h38f86fd4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c0; din <= 32'he6aa6989;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h126; din <= 32'he73f81be;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e5; din <= 32'hdb155b5c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h293; din <= 32'ha74d30fb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34d; din <= 32'hbbd15269;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h203; din <= 32'h3dbbbe8a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h178; din <= 32'h48c28282;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h070; din <= 32'hc300f51f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d9; din <= 32'h887aa9c5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h266; din <= 32'hc09eaa9c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h018; din <= 32'h9d27ce36;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e5; din <= 32'h6ce683e9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h016; din <= 32'h2506ba05;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h395; din <= 32'h314a45d5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f0; din <= 32'hb1715135;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h352; din <= 32'h9901b058;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b4; din <= 32'hf089468f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f5; din <= 32'h3996f382;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d8; din <= 32'ha4540c99;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h016; din <= 32'he6c3a95e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0dc; din <= 32'h689fc337;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04a; din <= 32'hfe5c9c3b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02c; din <= 32'h4305141d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03f; din <= 32'hd844a753;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15f; din <= 32'h18751ae9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e6; din <= 32'ha7b20fb5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b2; din <= 32'h79ba405c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33c; din <= 32'h4ab8e15f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b5; din <= 32'h50d36cbc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39d; din <= 32'hbd03e110;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d7; din <= 32'h2c476079;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h159; din <= 32'h20778fdc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18f; din <= 32'h61b43c9e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h239; din <= 32'h51c557c9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20e; din <= 32'h168aa688;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e1; din <= 32'h4c881f85;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h168; din <= 32'hfca36eef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d9; din <= 32'hfcc58c41;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a7; din <= 32'h7cc42547;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38f; din <= 32'hb105c358;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h366; din <= 32'h58a954db;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h339; din <= 32'he9e02705;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24b; din <= 32'hf9fa77e7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h064; din <= 32'h8e57f016;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e7; din <= 32'hdbd675cf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h299; din <= 32'h3e7f42f1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ff; din <= 32'hb9e4c10a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01d; din <= 32'hddbc7de9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33b; din <= 32'h7a377ac0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h343; din <= 32'h379704b2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h111; din <= 32'h7273ef02;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bd; din <= 32'h5af78576;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b4; din <= 32'hd78a1487;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15f; din <= 32'h601be067;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10e; din <= 32'h496933a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h201; din <= 32'h23d2bfcd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c4; din <= 32'h24f37771;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24e; din <= 32'hb25f7e5a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d8; din <= 32'h2a4c9f76;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13b; din <= 32'he6cff8ff;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07d; din <= 32'hba599cf2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0dc; din <= 32'h31560fa3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h269; din <= 32'hde5a929e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2df; din <= 32'h37583721;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f8; din <= 32'hd6d8cf5c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bf; din <= 32'hbc3d3f99;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e1; din <= 32'h65a28bac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h281; din <= 32'ha1440710;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h352; din <= 32'h2c281bbe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b4; din <= 32'he471db99;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e8; din <= 32'hf3147f9d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e3; din <= 32'h49aead2f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16b; din <= 32'h1b44286b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h330; din <= 32'h3b9efcc5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29c; din <= 32'h20bf4d04;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13f; din <= 32'h6b0109f4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h177; din <= 32'ha7c90dc0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a8; din <= 32'h61922650;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09a; din <= 32'hc22cd151;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h397; din <= 32'hfcceccf7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h087; din <= 32'ha3867862;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00b; din <= 32'h85db15eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17f; din <= 32'h0f8402ac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h304; din <= 32'h3fad15e2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bf; din <= 32'h9bb50068;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31c; din <= 32'hcb973456;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h393; din <= 32'hf53d226f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h019; din <= 32'hf902a594;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h396; din <= 32'h365de7bc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e7; din <= 32'h6685e12f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a0; din <= 32'he32d432d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a5; din <= 32'h73899f34;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h107; din <= 32'h6b5ba412;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36a; din <= 32'hc7ec693c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h234; din <= 32'h33dd3ca2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h287; din <= 32'h0f7087fe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h322; din <= 32'hd851bacb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d4; din <= 32'h4118338e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b8; din <= 32'h1f358118;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h200; din <= 32'h6bf956cb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e6; din <= 32'hdfdde551;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11f; din <= 32'h1168673c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d6; din <= 32'hdcbbb45a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3df; din <= 32'h6b644c6e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31f; din <= 32'ha2fbd5b1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39b; din <= 32'h199b003d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02e; din <= 32'h9a94fecd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2aa; din <= 32'h8a0e5796;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1da; din <= 32'h1561a50a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a1; din <= 32'h7081f2cd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c5; din <= 32'h8b315a3f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h067; din <= 32'haed9a708;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05e; din <= 32'h86f2a6f1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h350; din <= 32'h6cdc7a8a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h253; din <= 32'h15c60b32;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d5; din <= 32'h145d94d3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ce; din <= 32'h1cc1ba48;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ae; din <= 32'h7de46eac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h189; din <= 32'hac7051bf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30b; din <= 32'h88afce02;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h137; din <= 32'ha5e6403e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37b; din <= 32'h38738cd9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d8; din <= 32'ha08208e5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06e; din <= 32'hf1b8f9fb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h024; din <= 32'hc5c8ec97;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h207; din <= 32'h37ab7da7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31e; din <= 32'h9b81ff79;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h126; din <= 32'h7b388a79;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36e; din <= 32'hbde8687d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a7; din <= 32'h186f30d6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06d; din <= 32'hb0f1578e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h061; din <= 32'h5d99d260;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ee; din <= 32'h4de1e4b8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ce; din <= 32'h6ae2941f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d4; din <= 32'haceafe60;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cc; din <= 32'hca190ff9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05e; din <= 32'h393da539;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d3; din <= 32'h20dd50d6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d2; din <= 32'hd9569139;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d3; din <= 32'h58a5cb6d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h078; din <= 32'hc8a45a2a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h388; din <= 32'ha5881e87;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39f; din <= 32'h82aac544;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12f; din <= 32'h98564e27;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h143; din <= 32'hbe47d498;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07e; din <= 32'hcf6d6817;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h172; din <= 32'hb5e0c034;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b4; din <= 32'h5b871720;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h105; din <= 32'hce404656;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18b; din <= 32'h9b0b05bd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f0; din <= 32'h2569130c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e7; din <= 32'h53d3771a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0be; din <= 32'h6ef05732;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13d; din <= 32'h8a744076;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h143; din <= 32'h13c094af;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h220; din <= 32'haf730d1f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h228; din <= 32'hd2c4de3a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29e; din <= 32'hd0fef971;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h379; din <= 32'hd785032c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24c; din <= 32'h26170277;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h241; din <= 32'h48dfa50e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h195; din <= 32'h48f6dbad;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17c; din <= 32'h2b966a6d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h316; din <= 32'h9fc4d7d7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h228; din <= 32'hd5ef43eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h303; din <= 32'hd457f47c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d7; din <= 32'hf01a85f5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h301; din <= 32'heabe0563;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h033; din <= 32'he93bfa28;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ca; din <= 32'h7e3225e0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h038; din <= 32'hd6a14af8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f7; din <= 32'hfa694bf6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h208; din <= 32'hd816ca66;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21d; din <= 32'h90c2863a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b0; din <= 32'h532be1c9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h262; din <= 32'hbd74b201;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h223; din <= 32'hd1007c75;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h136; din <= 32'h353dd8be;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b5; din <= 32'hf9a7c5e4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17a; din <= 32'h052c4162;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a3; din <= 32'h6ba4abc0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ad; din <= 32'h8ec33f72;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17c; din <= 32'h84b0b340;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h228; din <= 32'hb26bce8d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24b; din <= 32'heb71eed2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11a; din <= 32'h20511613;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13a; din <= 32'hc3377cc3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h131; din <= 32'h537b145f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27e; din <= 32'hc1a4eeed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h259; din <= 32'hc83e2af3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c7; din <= 32'hf14b88cc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h393; din <= 32'h48172abd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c2; din <= 32'h71ead029;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01a; din <= 32'h24b3ba2a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c0; din <= 32'h2a2281f3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h173; din <= 32'heac8a345;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13a; din <= 32'h957e31dc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39d; din <= 32'hb0a7eb2e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31d; din <= 32'h11761a24;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f5; din <= 32'hf77cf129;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h178; din <= 32'h2d6131a3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h280; din <= 32'h7c0acbaa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a7; din <= 32'h2acadda6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26c; din <= 32'hb356fe7c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e4; din <= 32'h9df239ca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h039; din <= 32'h6e81ee92;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h243; din <= 32'h22f0389b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e7; din <= 32'h92a4985c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c0; din <= 32'h397deb56;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ac; din <= 32'h856211b0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h125; din <= 32'h7ecef011;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h169; din <= 32'h3fdba30a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h173; din <= 32'h89b94307;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h356; din <= 32'hf64fa617;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2da; din <= 32'hc0b9e958;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24e; din <= 32'hb10afda1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h178; din <= 32'h6aa0666f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h314; din <= 32'h3553ed8f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h310; din <= 32'hcb058321;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d7; din <= 32'h03264cff;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ce; din <= 32'h1e63b394;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h329; din <= 32'h93f0cfdf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30d; din <= 32'hbb32c84e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a0; din <= 32'heeae0757;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1dc; din <= 32'h33c790a4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fe; din <= 32'hcf9c18f1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09d; din <= 32'hffb855f6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h384; din <= 32'hb61110c7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09d; din <= 32'hb931649f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04d; din <= 32'hd7bf2c8c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b2; din <= 32'h8ba66d2f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ad; din <= 32'h03d59198;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h031; din <= 32'hb922bfbb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26c; din <= 32'h9b8d7f78;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33f; din <= 32'h32391a0f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d4; din <= 32'ha9c82ed3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29e; din <= 32'hebb34f7e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b8; din <= 32'h1b8b0323;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26d; din <= 32'h7df7c252;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h210; din <= 32'h6b1ba7d7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ae; din <= 32'ha3dfefdb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h389; din <= 32'ha0633c2d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37c; din <= 32'h16ade48b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28b; din <= 32'h760e2d09;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2db; din <= 32'h95c9b718;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h335; din <= 32'h3b105691;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h111; din <= 32'hcab0e638;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bd; din <= 32'hbd1759d2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a6; din <= 32'h170883c2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h053; din <= 32'hcab77f6f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00b; din <= 32'h53c114b9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h262; din <= 32'h1c940c4e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ff; din <= 32'h4eadc9d9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h085; din <= 32'h68b165a2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33b; din <= 32'ha6092058;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f1; din <= 32'h86a60de9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33b; din <= 32'hc3312e5d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d8; din <= 32'h268de35c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h139; din <= 32'hc79f013a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34f; din <= 32'h857afc5e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e2; din <= 32'h6c969411;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2fd; din <= 32'hd9666025;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h283; din <= 32'h784616bd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d3; din <= 32'hda95e7b2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3de; din <= 32'hc97bd880;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h156; din <= 32'hbb799e2e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h274; din <= 32'hd66baf6e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h081; din <= 32'hf78af22e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b6; din <= 32'h32525325;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06f; din <= 32'h54c2a19f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h317; din <= 32'h5482d289;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ae; din <= 32'h5b43c19f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04a; din <= 32'h4c80565a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3df; din <= 32'h05ee02ef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h354; din <= 32'h7c476d44;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b4; din <= 32'ha0da282d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16d; din <= 32'hf65f443e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h000; din <= 32'hcc24477d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h022; din <= 32'hf2eb31aa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e2; din <= 32'h7cfe43d6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h154; din <= 32'h67c6ec4b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36f; din <= 32'h6087e771;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31e; din <= 32'hb492b150;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09c; din <= 32'h57bfffd9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b9; din <= 32'ha53cef80;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h099; din <= 32'hf0b51a15;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h252; din <= 32'hfa35bc2c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12c; din <= 32'h255194c9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cf; din <= 32'h4d305aec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h355; din <= 32'h13ca2c4a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38d; din <= 32'h125f885b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h338; din <= 32'h3011a8bf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12d; din <= 32'h2049cde0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0aa; din <= 32'h8da5e618;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h133; din <= 32'h5dfd9df8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fa; din <= 32'hf8577d21;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a9; din <= 32'h5bf087c5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h251; din <= 32'hd374d0fb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h211; din <= 32'hf9e2a6b1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h278; din <= 32'hc731aa4b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f4; din <= 32'h1fe07976;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h282; din <= 32'hf13149c6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20c; din <= 32'h0583f5a1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h359; din <= 32'h13eca0fe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29e; din <= 32'h3d6ae636;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39f; din <= 32'h646d66d2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h142; din <= 32'hd9201e53;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fa; din <= 32'h1f237b0a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ad; din <= 32'hb1eb7f95;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h167; din <= 32'h42c7690e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h347; din <= 32'hdabbb99b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h118; din <= 32'h9b9d40e9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e3; din <= 32'hda9d4efb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h305; din <= 32'hf8caf533;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c2; din <= 32'h7a6f140d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h067; din <= 32'h2a773d65;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h051; din <= 32'hd9e5bf88;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h181; din <= 32'hfc0482d1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a8; din <= 32'h40082afb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f1; din <= 32'h0c487021;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26f; din <= 32'hf96d01d2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a8; din <= 32'h7575c785;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h034; din <= 32'hc9472c88;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h206; din <= 32'h407477c1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29a; din <= 32'h73d9c8d4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09b; din <= 32'h420a03da;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h338; din <= 32'h2e9679d9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h373; din <= 32'ha93ae8f5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h002; din <= 32'h5e989bcb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h385; din <= 32'hab57b3d3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3dd; din <= 32'heb9069e4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c2; din <= 32'h66b511ed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12d; din <= 32'h5fe6f41d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f6; din <= 32'h8dd9a4fc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d3; din <= 32'h132eb211;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13d; din <= 32'h714b4a4c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d9; din <= 32'h60cae29c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h239; din <= 32'h6c0d43d2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22e; din <= 32'h0ff41f2f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h239; din <= 32'h1b5aef4e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a1; din <= 32'hdbf2bc95;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h398; din <= 32'h0942bc6c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h303; din <= 32'h0b17b426;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fd; din <= 32'h78ddda75;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h011; din <= 32'h392e39b6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ff; din <= 32'h8285443a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h228; din <= 32'h2f7c0d8d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26f; din <= 32'hcc440b73;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e2; din <= 32'hf98bde7f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h134; din <= 32'hc4e85215;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h327; din <= 32'hde144ff9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22c; din <= 32'h1f06d048;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b5; din <= 32'h48ef937c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02b; din <= 32'h9356ea08;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a9; din <= 32'ha76df8f9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ef; din <= 32'h09433c2a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h119; din <= 32'h05b1b7e4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h254; din <= 32'hf782294f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e0; din <= 32'hc78ec9cf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h266; din <= 32'h33d5e318;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0be; din <= 32'ha9144889;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h186; din <= 32'h7af0a2c1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b4; din <= 32'h4795af0e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e7; din <= 32'hd5fe9a7a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b0; din <= 32'h00b914a2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bc; din <= 32'h9d433f21;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h128; din <= 32'h42c8fd91;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d7; din <= 32'hfd75c14a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h304; din <= 32'h4cc0ccab;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04c; din <= 32'h4a48effc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h390; din <= 32'h7dc27106;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12f; din <= 32'h319a3400;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h239; din <= 32'h077eaacc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29a; din <= 32'h264babde;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24b; din <= 32'hb8ab39fd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h208; din <= 32'h2435c66c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c2; din <= 32'hf70899bd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35d; din <= 32'h9ebd8c72;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h128; din <= 32'h400c81b1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h158; din <= 32'hb930ad3b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h092; din <= 32'h45c0f201;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d1; din <= 32'h94e21a58;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h348; din <= 32'h675c50aa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cd; din <= 32'hdd6b6755;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h107; din <= 32'hd172dba3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e0; din <= 32'h0d080b1a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h054; din <= 32'h7888b539;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h082; din <= 32'h051205df;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37c; din <= 32'h2e9349d0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22e; din <= 32'hf9c6a630;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f1; din <= 32'he9ab4319;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10b; din <= 32'h0c792442;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h098; din <= 32'he2fcd2b7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33c; din <= 32'hbe072537;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07f; din <= 32'h8eca868e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d7; din <= 32'h6364f675;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h007; din <= 32'h060ce05e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c4; din <= 32'h0b57be11;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11e; din <= 32'hc0836665;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h122; din <= 32'h50d86dc4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ba; din <= 32'hb99175f5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h185; din <= 32'h730735e9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e8; din <= 32'h7c8b2938;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h239; din <= 32'hbd3b2e24;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39c; din <= 32'h50e406d0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h267; din <= 32'hc0026ea7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35c; din <= 32'h1fbda2d3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h023; din <= 32'h3c93ed42;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h333; din <= 32'hf2b8bad7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h049; din <= 32'hbaf26c9b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h330; din <= 32'h274bfb19;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bf; din <= 32'hf8b43e8c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31e; din <= 32'h7820c246;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a2; din <= 32'h3ae4bac0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a4; din <= 32'h958ba15d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h391; din <= 32'hfcffa4fe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ed; din <= 32'h8cb35849;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24b; din <= 32'h6d35275e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h320; din <= 32'h4e46adea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c1; din <= 32'h1ff96832;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1db; din <= 32'ha923c94c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c0; din <= 32'h83108ccb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h179; din <= 32'h654edb57;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3af; din <= 32'hdc9a251f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f3; din <= 32'h4bb456d8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f5; din <= 32'ha8a3b87d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35a; din <= 32'hb49b1b09;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h241; din <= 32'hb8827fdf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h382; din <= 32'hcad1e20a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c3; din <= 32'ha1373b88;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ef; din <= 32'hc3828461;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h247; din <= 32'h66a33fd3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3df; din <= 32'h67e04a46;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h245; din <= 32'h217b2981;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h226; din <= 32'hbd26e9dc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h131; din <= 32'h39feabd6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h155; din <= 32'hb0c4a53f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b0; din <= 32'h570574af;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fe; din <= 32'h28efd4d4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h300; din <= 32'h8aaf374c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3da; din <= 32'h9cde75ee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b3; din <= 32'hc3029404;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cf; din <= 32'h7aaf9c76;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cc; din <= 32'h74c85506;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h381; din <= 32'h5b8fcd51;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38c; din <= 32'hd2f1d21c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h083; din <= 32'hacff5447;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h266; din <= 32'hcb551acd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e2; din <= 32'h162c275c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h096; din <= 32'h1d8e618e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a4; din <= 32'h91dba65f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c6; din <= 32'h3abe53f7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08d; din <= 32'h782868bf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h003; din <= 32'h37bd3012;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h167; din <= 32'h92a7a537;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34c; din <= 32'h3dc3af7d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h086; din <= 32'hfc6bfe3e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30f; din <= 32'hf279bc13;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h300; din <= 32'hd95b4caf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h107; din <= 32'hfd587425;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29d; din <= 32'hd40a6e9e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06d; din <= 32'hb81f6a55;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06a; din <= 32'h8bdd163d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h021; din <= 32'h3511cca3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h113; din <= 32'h10a88b83;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ad; din <= 32'h68eb2d2b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f9; din <= 32'h7929bafc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a0; din <= 32'ha9e27f50;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h270; din <= 32'h27c5579b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00c; din <= 32'h7b86c9f4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h367; din <= 32'h70fe3d5e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e0; din <= 32'h96325f32;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a0; din <= 32'h5f249dfc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07f; din <= 32'hfa47637d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h062; din <= 32'h7ecaeb03;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d4; din <= 32'h17d40b31;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h166; din <= 32'hbc1c4cbe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d7; din <= 32'hbc484635;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10f; din <= 32'h1dee3437;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1da; din <= 32'h2bb55bf9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a8; din <= 32'he2091aec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a9; din <= 32'h89adc83b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a9; din <= 32'h51fc3686;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h054; din <= 32'h861e165d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h034; din <= 32'h11c3a466;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15e; din <= 32'h9d1f4485;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a8; din <= 32'hf6573672;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h219; din <= 32'h91e7741e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a0; din <= 32'h19cc1f91;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h031; din <= 32'hdba46c35;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36e; din <= 32'hb83f66fa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bc; din <= 32'hd43b3d71;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20a; din <= 32'h534c3bef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h182; din <= 32'hfe846c13;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b8; din <= 32'h426f1ae2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03f; din <= 32'h6c0cd3a1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b3; din <= 32'h85b7f001;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16c; din <= 32'h687c5261;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h107; din <= 32'h09215224;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h137; din <= 32'hc99794a8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a4; din <= 32'h6a3fb6ef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a8; din <= 32'hcd5f9901;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a5; din <= 32'h1dbb1208;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h218; din <= 32'h5723ffd7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b3; din <= 32'h7c789e54;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h061; din <= 32'h9e432457;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h278; din <= 32'h4b8fef9b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h152; din <= 32'h5aa917aa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d1; din <= 32'h833d27c3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h171; din <= 32'h552b12f7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b4; din <= 32'haaa408a1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fe; din <= 32'hc18e899c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05d; din <= 32'h01ea7187;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ea; din <= 32'h640c1ea6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25d; din <= 32'h1a37c0a7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39f; din <= 32'h69148435;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h050; din <= 32'hc3469b3e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h293; din <= 32'h3f19ecba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c9; din <= 32'h6daf3118;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b3; din <= 32'he4850071;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39a; din <= 32'hec088d1e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37d; din <= 32'h4c0295c5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h252; din <= 32'hc3e93abd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f2; din <= 32'h5c3ef462;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b1; din <= 32'ha4aae182;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ad; din <= 32'h4e325088;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a6; din <= 32'hbbd9f255;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ef; din <= 32'hcbf70530;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ad; din <= 32'h615c1744;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11c; din <= 32'ha770e883;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00d; din <= 32'hdf87e92f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ea; din <= 32'h21ac7f7f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h209; din <= 32'h8d894075;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b8; din <= 32'h5739b648;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h306; din <= 32'hcc82df0b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39f; din <= 32'h88457823;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b4; din <= 32'h935dbba5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bd; din <= 32'hb2aac1fb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h396; din <= 32'h48110ebe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ca; din <= 32'hcf13474b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00f; din <= 32'hfc5ade2e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b4; din <= 32'hff9d131d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bf; din <= 32'hfb4f533b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ea; din <= 32'h46192928;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30b; din <= 32'he09cebd4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h236; din <= 32'h9b7d7800;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d5; din <= 32'h6c7007d6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32d; din <= 32'hc0f6e7e1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09e; din <= 32'h37861e53;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h335; din <= 32'hd50689e8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d4; din <= 32'h6ec4060d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h095; din <= 32'hfecfe8cf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cf; din <= 32'h481f3103;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d2; din <= 32'h3a12ed4a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d9; din <= 32'h734722ed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18a; din <= 32'hc66f366f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a1; din <= 32'hee8f5520;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b7; din <= 32'ha5bdd6b9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08a; din <= 32'h288302cb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h249; din <= 32'hd1e18c56;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h092; din <= 32'h5124bf84;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03b; din <= 32'hfed985e5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h398; din <= 32'he0d85d1b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14c; din <= 32'h046e1136;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39a; din <= 32'hc0217ab2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2dc; din <= 32'h18297568;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32f; din <= 32'h1bd2a57e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cb; din <= 32'hdcb75b6c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ef; din <= 32'h7a93bfd4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h137; din <= 32'hd3f9ef4b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1eb; din <= 32'h81c46eb7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cc; din <= 32'hf037a202;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b2; din <= 32'hfd89d3f5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d3; din <= 32'hf64e8ed2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h366; din <= 32'h2042c1ab;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37e; din <= 32'h26b74e02;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30b; din <= 32'h754fd2de;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h305; din <= 32'hb191a0eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37a; din <= 32'h0ec38532;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h323; din <= 32'h63ee57ec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bd; din <= 32'h3f704a65;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h354; din <= 32'h8020fa53;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1db; din <= 32'hda167d76;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15b; din <= 32'h07c37887;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bf; din <= 32'h372a5878;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b8; din <= 32'hcb0f598a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h139; din <= 32'h04b59ba2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h134; din <= 32'hb2bc5b69;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b4; din <= 32'h8300ef05;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a5; din <= 32'h4ae88213;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cf; din <= 32'hc351b24b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h314; din <= 32'h53f303b9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07b; din <= 32'he5e24644;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h156; din <= 32'he1a2e3b2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h253; din <= 32'h30010499;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d1; din <= 32'hc56e92d2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h186; din <= 32'h2ad64f63;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a3; din <= 32'hc603bc06;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h073; din <= 32'haffcb9c7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ea; din <= 32'hbfe67e4a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h267; din <= 32'h0d18f046;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h335; din <= 32'h7bbbe312;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h370; din <= 32'h66d57ae6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h045; din <= 32'he1f4c1ca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a9; din <= 32'hf1d1531f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a8; din <= 32'hd46293e7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h204; din <= 32'h1121196b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ee; din <= 32'he742a48d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h077; din <= 32'h636a924d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02c; din <= 32'h075cbf01;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03a; din <= 32'h9dca5a8a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15a; din <= 32'h5600d24e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c2; din <= 32'hfe6ad47d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h167; din <= 32'h572c16ab;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h373; din <= 32'h6cafc382;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e1; din <= 32'ha1552a9b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cf; din <= 32'h58c8121a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h148; din <= 32'hc1d9b1bd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f6; din <= 32'h3fa33d21;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h050; din <= 32'ha0c3cabd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b7; din <= 32'hceada374;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22f; din <= 32'h0fd5c1f8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h291; din <= 32'h5b186b37;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cf; din <= 32'h57f97227;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h380; din <= 32'h7a65047f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38f; din <= 32'h116c3572;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h018; din <= 32'h5aa9cb86;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c5; din <= 32'h9ac509ca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d4; din <= 32'hdeea6ae4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h126; din <= 32'h24190424;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h311; din <= 32'hc380db58;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a6; din <= 32'h8b608ef0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b1; din <= 32'he5c10703;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h277; din <= 32'h69f318b7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h069; din <= 32'hca6a1dbc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29d; din <= 32'h14829d8c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ce; din <= 32'h291d6ee0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c2; din <= 32'h544727b7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20a; din <= 32'he554ea66;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0aa; din <= 32'hb065dfca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b7; din <= 32'he04ec954;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h190; din <= 32'h94c5824d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cf; din <= 32'ha7f4e971;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c1; din <= 32'h43abec4a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h132; din <= 32'h2e3a6b80;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a5; din <= 32'h82ea55ed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17a; din <= 32'h8496aa79;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h337; din <= 32'h3f69c8ac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c1; din <= 32'h78845e89;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f4; din <= 32'h068c22ba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a5; din <= 32'he79a6b35;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26f; din <= 32'hbdb178e4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10e; din <= 32'hb02eb508;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b1; din <= 32'h4abb38fb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h279; din <= 32'h2fdbc8ae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h055; din <= 32'ha115fc09;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b4; din <= 32'he283f865;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3df; din <= 32'h17cdd6d7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ea; din <= 32'hd9edbed4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cf; din <= 32'h781aee5d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h222; din <= 32'h5c7e1fd0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c4; din <= 32'h4128147d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d5; din <= 32'hbdd20658;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h226; din <= 32'hdfbed817;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38d; din <= 32'h8ec5a470;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h081; din <= 32'h39a6eb83;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h350; din <= 32'h423db497;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33f; din <= 32'hb618d75d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h078; din <= 32'h919b3c7b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h112; din <= 32'ha4f4cef4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15d; din <= 32'he2732851;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h034; din <= 32'he2e2e46c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d2; din <= 32'hbdf3f3ee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e3; din <= 32'h97ac626d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b4; din <= 32'h2b839916;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h010; din <= 32'h7f033417;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f3; din <= 32'h1243abbc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03a; din <= 32'h127d4461;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h053; din <= 32'hc100b5fd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23c; din <= 32'h6e6f89e5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h291; din <= 32'h82504338;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20d; din <= 32'h4d026a1e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25f; din <= 32'ha19cc70e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h070; din <= 32'hfb3346f5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0be; din <= 32'h1bf92a61;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h039; din <= 32'h8c63171a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h077; din <= 32'hbf8ca4b2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f0; din <= 32'hf8a3bfe1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bd; din <= 32'h29d94f6d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22d; din <= 32'h71f4b7a8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c8; din <= 32'ha3959f38;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h196; din <= 32'h66140ced;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h385; din <= 32'h41bd4db8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h316; din <= 32'h0905ed6a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e6; din <= 32'h683363d2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h007; din <= 32'hfbf85ef8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h259; din <= 32'h5db8d6df;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a3; din <= 32'h8fe071d7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ed; din <= 32'hed57e448;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f5; din <= 32'h0cfaae78;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02b; din <= 32'hf926f469;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h334; din <= 32'hb916d307;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h045; din <= 32'hae18448b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27c; din <= 32'h813c95c3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h239; din <= 32'h9966905f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09e; din <= 32'h4105f0f7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h052; din <= 32'h34387663;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h084; din <= 32'hb4a864d8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h099; din <= 32'h68cd5675;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h387; din <= 32'hd5386533;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ed; din <= 32'h3beb3c92;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h178; din <= 32'h33eecbbe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h256; din <= 32'h5ca4fbd3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h276; din <= 32'ha7d41a9d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f3; din <= 32'hb5ba4789;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d0; din <= 32'hb128f765;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06a; din <= 32'h0ac7d45b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h152; din <= 32'hf18f2256;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13d; din <= 32'hb8ad7247;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h349; din <= 32'h141e96d4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d9; din <= 32'hbd18e188;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e5; din <= 32'h36fb7f60;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h233; din <= 32'h86062e7d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h112; din <= 32'h4d4a913a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h194; din <= 32'h3778585e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17b; din <= 32'hc2d7d639;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b0; din <= 32'h831f44ba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ab; din <= 32'hcf072132;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cf; din <= 32'he96f4c6e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h156; din <= 32'hca83be4b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h115; din <= 32'hf43b234e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d5; din <= 32'h5e70c1ba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19c; din <= 32'he0b64d81;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h181; din <= 32'h32559b18;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h277; din <= 32'h1efe840c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37c; din <= 32'hf2fae77b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h255; din <= 32'h1a25835a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h298; din <= 32'hb5d3433b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24b; din <= 32'h6dc882c1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15f; din <= 32'hb6e3c71b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ed; din <= 32'h994d54f9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f5; din <= 32'hedba5605;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f0; din <= 32'hdaf5c413;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h345; din <= 32'h1aff47c2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24d; din <= 32'h3bd81e96;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a5; din <= 32'hab41640c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h106; din <= 32'h79666606;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h267; din <= 32'hbe82066b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fb; din <= 32'h9be88d5a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d0; din <= 32'hfe7ac7a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09d; din <= 32'hdff0770c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11a; din <= 32'hd265a285;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15a; din <= 32'ha4aa43a7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h157; din <= 32'h1b7ed1ee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f1; din <= 32'h7b2f49d3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11a; din <= 32'h9b8168f1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c7; din <= 32'h4e9c5e28;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d3; din <= 32'hb7faafca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h378; din <= 32'h78d62220;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21c; din <= 32'heee51bc7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h362; din <= 32'h72f84540;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c6; din <= 32'h90ad0b49;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19f; din <= 32'hd228aaa8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d7; din <= 32'he308b1ec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h330; din <= 32'h4c968a96;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h326; din <= 32'h06ecab7c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a8; din <= 32'h0ccc5059;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h029; din <= 32'hcd86d342;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3de; din <= 32'h95a9e879;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24e; din <= 32'hbc7f4623;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22f; din <= 32'hd9d481e7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33e; din <= 32'hcc8f19d4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f8; din <= 32'h1d75ca9a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h343; din <= 32'hef3ef2e2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a1; din <= 32'h38726bc2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h153; din <= 32'h211a263a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h087; din <= 32'h89d8e21f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a0; din <= 32'hd72f18a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ca; din <= 32'hb080522d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h344; din <= 32'hafc6b394;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a6; din <= 32'h4a41788e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15a; din <= 32'h506982cd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16b; din <= 32'hdd342bfc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c6; din <= 32'he5fd57c0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h089; din <= 32'hdebc3246;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36e; din <= 32'h416df8cf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e8; din <= 32'h32120342;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16d; din <= 32'h15f63e39;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h065; din <= 32'h84609518;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04b; din <= 32'h7ea12003;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h123; din <= 32'h31023deb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e2; din <= 32'hc3d27ddd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03f; din <= 32'h74e9a06a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e6; din <= 32'hcec9f826;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2fc; din <= 32'hd95147b8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bc; din <= 32'h0de9cc92;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h016; din <= 32'h4f1ba318;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h285; din <= 32'h8304605a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h056; din <= 32'h14cdf88f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h364; din <= 32'hea53ae60;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a4; din <= 32'he0cfebf0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32e; din <= 32'h2081aed7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h200; din <= 32'h15bacce2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h039; din <= 32'h625266bc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b5; din <= 32'ha128fe1f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h047; din <= 32'hc00aa302;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32f; din <= 32'h6362136d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h247; din <= 32'h7d7c6815;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ea; din <= 32'hb02d5bd5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h151; din <= 32'h94a00344;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h389; din <= 32'h8362cd24;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ec; din <= 32'ha4283d63;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00a; din <= 32'h93fa8020;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09a; din <= 32'h5ec5ac4e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1df; din <= 32'h7c06d5fd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h009; din <= 32'haa1c735a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cd; din <= 32'h237e80e7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h364; din <= 32'h9b249631;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h052; din <= 32'hde6b3718;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h161; din <= 32'h63c309e8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fa; din <= 32'h2669b79b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b2; din <= 32'h11111603;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h074; din <= 32'hd9e72d27;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32a; din <= 32'h17a14cee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h347; din <= 32'hfe1f2f91;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h351; din <= 32'h82109184;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d2; din <= 32'h20a041f7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32f; din <= 32'h81735c3b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h204; din <= 32'hb146ce09;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b3; din <= 32'hea25ac0e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d3; din <= 32'h090781f6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h198; din <= 32'h3290c6f6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h161; din <= 32'hf7175906;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a0; din <= 32'h92c06ab8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39f; din <= 32'h521d4c1b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h383; din <= 32'h7abbde6b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22e; din <= 32'hbc79be70;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h231; din <= 32'haedd2cd9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b1; din <= 32'h9bde60e6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h190; din <= 32'hcfab28ff;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07d; din <= 32'h306f539b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fb; din <= 32'h8fb291b9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h232; din <= 32'he04b8963;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h096; din <= 32'he82a91e2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23e; din <= 32'h65dfbcf6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h039; din <= 32'h4207c99d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1eb; din <= 32'he847c7ab;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h098; din <= 32'he03bdbb0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bf; din <= 32'h9b52e93c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f0; din <= 32'he868c428;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h061; din <= 32'h8699ed2a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a6; din <= 32'h7024d53a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09e; din <= 32'h0e10c0ac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ee; din <= 32'h7d4db79a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07f; din <= 32'h0697d7ff;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fe; din <= 32'h1919a8e2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h012; din <= 32'h1f7edf14;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a5; din <= 32'h000ff08e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h039; din <= 32'haad8a8e4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h282; din <= 32'h724984a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bb; din <= 32'hd0a1f293;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c4; din <= 32'hebb307d5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22b; din <= 32'h19d452ef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37e; din <= 32'h6391c87a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h204; din <= 32'h7da8d4ca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bc; din <= 32'hec0b3b11;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b1; din <= 32'h1144f0d9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38b; din <= 32'h113ed768;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h381; din <= 32'h12b39c3c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e5; din <= 32'h431dc1ef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2db; din <= 32'ha2e53227;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12f; din <= 32'h0c7b092f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b5; din <= 32'h1085a458;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h244; din <= 32'h3c2c92cd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2fb; din <= 32'h9f9722e0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36f; din <= 32'h704d6ec8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h366; din <= 32'h5a31547c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h106; din <= 32'h982691dd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14e; din <= 32'hacfc5110;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e4; din <= 32'h0a62291f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a0; din <= 32'hb2eb1ac1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h296; din <= 32'h531dd482;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a7; din <= 32'h855c368c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e2; din <= 32'h060648f2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07c; din <= 32'h9f551882;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07c; din <= 32'hda5976e4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ee; din <= 32'hc095e19b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h359; din <= 32'h75b1053d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h289; din <= 32'h6145637b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a7; din <= 32'h4cf3a9f6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d8; din <= 32'h4b7f1405;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h384; din <= 32'hf5a4dcec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h342; din <= 32'ha1334484;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38f; din <= 32'hf1d41ef0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h039; din <= 32'h78e579b9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h059; din <= 32'hddd4731b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c2; din <= 32'h63ea8d90;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a5; din <= 32'h8812ec80;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2da; din <= 32'hc64537a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29a; din <= 32'h327fe830;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h374; din <= 32'h78746c44;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d2; din <= 32'h0bace6ad;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36d; din <= 32'h864af206;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36b; din <= 32'hc5124c2f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h317; din <= 32'h927ef405;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09e; din <= 32'h45356be2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24f; din <= 32'hfc354cd3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d4; din <= 32'h25fe7e83;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h033; din <= 32'hbef6e9be;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ea; din <= 32'hd3bebc70;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h216; din <= 32'h89f1874a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h026; din <= 32'h1cdc5a30;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h106; din <= 32'h8b88e8df;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18c; din <= 32'hd4cc5a48;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d8; din <= 32'hcd490e45;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h331; din <= 32'hd06f2361;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29f; din <= 32'h8a5b0b9b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23c; din <= 32'h9ded2d8a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3dc; din <= 32'h13809b02;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26e; din <= 32'hf1a06c65;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h139; din <= 32'h3db13bc0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cb; din <= 32'h7b62a3f6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h111; din <= 32'h7afc4457;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cd; din <= 32'hc18e76ea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h249; din <= 32'h9f319dee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2fa; din <= 32'h79ee0397;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a5; din <= 32'h253df8d9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h062; din <= 32'h9d6c0268;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ca; din <= 32'h2db59b9d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h079; din <= 32'h289cd92f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h265; din <= 32'h51c6c92b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d9; din <= 32'h5484f864;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e0; din <= 32'h99e98557;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b5; din <= 32'h593cd69d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34f; din <= 32'h6bab93f1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ff; din <= 32'ha401fe8f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27d; din <= 32'h88510bc8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c7; din <= 32'h33859f70;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h018; din <= 32'ha8bd9509;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f8; din <= 32'hd32a7371;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h193; din <= 32'h7d456385;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h140; din <= 32'hcde03ac3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13d; din <= 32'ha52ef5d4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0aa; din <= 32'h6de65afc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h354; din <= 32'h638a6295;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12d; din <= 32'h6c35280a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18e; din <= 32'h2bc21625;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c7; din <= 32'h3a3cbcfa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ce; din <= 32'h19dfc901;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e0; din <= 32'h03f6145d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h200; din <= 32'h433feaa4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e9; din <= 32'h8bc22d4e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34b; din <= 32'h9721907f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h333; din <= 32'hf3f1ebb2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34a; din <= 32'he842711f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h390; din <= 32'hb076a071;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h252; din <= 32'he307a300;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h297; din <= 32'h85894367;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h339; din <= 32'h511208f2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h249; din <= 32'hd3c6ad4e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h245; din <= 32'h7a31e52e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02e; din <= 32'h2ef0dfe2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h318; din <= 32'he200e8ea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h372; din <= 32'h71ca1704;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b2; din <= 32'h385e9f8b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h021; din <= 32'h10e2009f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h264; din <= 32'h77f67f17;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19a; din <= 32'hddfcd12b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h221; din <= 32'hffa6c19e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h257; din <= 32'h96dbd672;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25c; din <= 32'h304b3226;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b3; din <= 32'hc3deb8ec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29d; din <= 32'hae2bdf49;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c4; din <= 32'h5bf5d9af;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h140; din <= 32'h777a4d63;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h040; din <= 32'h8bcc00bb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27e; din <= 32'hf1d04683;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e5; din <= 32'h8afb2d62;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h291; din <= 32'h4283f2d9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2eb; din <= 32'hf739f482;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0df; din <= 32'ha2bebc20;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37f; din <= 32'h78b3faf0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28e; din <= 32'h8e5241db;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e8; din <= 32'h630c56e7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cc; din <= 32'h586a1c7f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h334; din <= 32'h1cb29c81;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h135; din <= 32'h69e0a30d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h151; din <= 32'h5196953c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ce; din <= 32'h95b84a2b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e0; din <= 32'h014554e8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h017; din <= 32'hca7675cc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a5; din <= 32'h5d8f17bc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d6; din <= 32'h33479001;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39b; din <= 32'hac46818b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ce; din <= 32'h5998ff5f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26a; din <= 32'h1c18b8e8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13b; din <= 32'h5d188434;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h159; din <= 32'h2c57d743;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h336; din <= 32'heada7585;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h016; din <= 32'h1e4684bc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h072; din <= 32'hc8f7dc3d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28c; din <= 32'h5921e01d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h189; din <= 32'hbb7b2a9b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h239; din <= 32'h67ba64a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f1; din <= 32'h1edd8fcf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23f; din <= 32'h84adc241;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20b; din <= 32'h21a32d00;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h286; din <= 32'h9d62d461;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ca; din <= 32'h137d03a4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ab; din <= 32'ha13b5a1b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b8; din <= 32'ha0a0d76f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h110; din <= 32'hda38954a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e9; din <= 32'haa5719de;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d8; din <= 32'h802f331c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h152; din <= 32'hc77d8107;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04b; din <= 32'hfc91a209;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25f; din <= 32'h97c87293;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h245; din <= 32'h9b16f97a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h093; din <= 32'hd8819a75;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2da; din <= 32'hb87f414f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a4; din <= 32'h29771470;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h279; din <= 32'hd6a33455;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c8; din <= 32'h83908733;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08f; din <= 32'h51c41088;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h240; din <= 32'ha5e09d7a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f9; din <= 32'h4f5bb14e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fb; din <= 32'h0978e0b4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28e; din <= 32'hd8de1b31;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h168; din <= 32'he7326b57;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d7; din <= 32'h7decac4c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f9; din <= 32'h99194d30;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h063; din <= 32'h1746a061;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03b; din <= 32'hb8bf553f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32d; din <= 32'h7ccf4d7d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h319; din <= 32'ha4b85e0e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h179; din <= 32'h0fab3ada;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h178; din <= 32'hb2659385;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27c; din <= 32'h3cba2be2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h281; din <= 32'h65bb6ff9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h210; din <= 32'hc1b3e087;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h242; din <= 32'ha8a1886f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a8; din <= 32'h2055f8df;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h141; din <= 32'h3100eddd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h011; din <= 32'h1f204622;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e1; din <= 32'h9cc73798;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d6; din <= 32'h6f123069;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c0; din <= 32'h50bacecf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h332; din <= 32'h424c83a3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h119; din <= 32'h8ba5d0d3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e4; din <= 32'h7f79d122;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17c; din <= 32'hafa9d978;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b5; din <= 32'h7bac2fe8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07d; din <= 32'h9f71ccd4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20f; din <= 32'h363d7ff7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h249; din <= 32'hba6dcac8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32d; din <= 32'ha681805e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h221; din <= 32'h5a26edc5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d6; din <= 32'hf7bc6a13;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0af; din <= 32'hb17ce62a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e9; din <= 32'h7322daec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ff; din <= 32'he8015299;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h380; din <= 32'h074af06d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26b; din <= 32'h1a2babcc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25e; din <= 32'h007af264;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h279; din <= 32'h29c09713;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25d; din <= 32'h969b726d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fb; din <= 32'h7e98a07a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h126; din <= 32'hdf88affe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e1; din <= 32'h0dd4ba53;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b8; din <= 32'h99b62ba1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h304; din <= 32'h442418c7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h065; din <= 32'h6e0764fb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h336; din <= 32'h5726eccf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d8; din <= 32'hae583aa6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h098; din <= 32'h6fe39199;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h345; din <= 32'h699d5db8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b5; din <= 32'h25b0c382;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h369; din <= 32'h122436b4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c7; din <= 32'h7b198d21;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h264; din <= 32'h62bc5f06;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10c; din <= 32'hc02658a3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ef; din <= 32'h9f034f13;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b1; din <= 32'h8ca6455e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a1; din <= 32'h274da93b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27e; din <= 32'hdf94e70f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h292; din <= 32'h285013c9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b8; din <= 32'h99981fb4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b9; din <= 32'hb220e4f6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e8; din <= 32'h0b2cc82e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09a; din <= 32'ha1462842;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h377; din <= 32'hdffa481c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h276; din <= 32'hc513f860;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ec; din <= 32'hf640fbc7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04b; din <= 32'h2589c81b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h057; din <= 32'h78b7c74b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bd; din <= 32'hdba84a88;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16a; din <= 32'h048d7014;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h191; din <= 32'h53287ae3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h271; din <= 32'h06139f7b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h272; din <= 32'h40655fe8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c4; din <= 32'he726d892;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b6; din <= 32'h0609f415;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27a; din <= 32'hc1f3d3dc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d5; din <= 32'h10aec6fd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h034; din <= 32'h2e686139;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h224; din <= 32'h9c8ce944;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38d; din <= 32'hfa2cb7f5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37b; din <= 32'h25f7366b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fd; din <= 32'h734dd92f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ff; din <= 32'h9a1fe3a3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h339; din <= 32'hc22d6a61;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f2; din <= 32'h656888f7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29c; din <= 32'h634e48cd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2aa; din <= 32'hc1a14b67;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h189; din <= 32'h24f4455a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h303; din <= 32'h4bfebb74;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f1; din <= 32'hf0813ca9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h003; din <= 32'h44b3df9e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h053; din <= 32'h4041b7a2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03d; din <= 32'h10a77f48;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d9; din <= 32'h7bd9d6b7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h192; din <= 32'h713ac39c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h360; din <= 32'h12caa472;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30d; din <= 32'h117c7406;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h171; din <= 32'h0e6237cb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22a; din <= 32'hfecf410c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2da; din <= 32'h309215f1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h350; din <= 32'h747299d0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h175; din <= 32'he51ae036;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13b; din <= 32'h033fd319;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fd; din <= 32'hfeda15e5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c5; din <= 32'h2c6c4a38;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21e; din <= 32'h85683487;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b4; din <= 32'hccedddcb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a0; din <= 32'ha39ba0e3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h383; din <= 32'hcf278180;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00f; din <= 32'h00e5f27c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h285; din <= 32'hbd7a8795;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0eb; din <= 32'h5a3e99fe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12e; din <= 32'h17d9481c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h117; din <= 32'h0986196e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e6; din <= 32'h52725c7b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17e; din <= 32'ha12d0ad1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fc; din <= 32'hf4157ab9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b0; din <= 32'ha3766fc4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f0; din <= 32'hb48425cf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h226; din <= 32'ha7a71066;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a6; din <= 32'h91dfbae9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31b; din <= 32'h664cbf4c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e6; din <= 32'h6c91a3f2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ed; din <= 32'h1e3037fe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h339; din <= 32'h99c92a93;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h257; din <= 32'h0aabcbde;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c7; din <= 32'h1bdf895e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h066; din <= 32'ha6c000c8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a0; din <= 32'h494b6829;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b9; din <= 32'h9ee44f9b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06c; din <= 32'h2af160a8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h146; din <= 32'h74fcac00;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h380; din <= 32'hb8d8deb4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3df; din <= 32'h18450766;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ca; din <= 32'hd8f48976;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1eb; din <= 32'hf8e14ba6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00a; din <= 32'h8cc1e7f4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23f; din <= 32'h3d4a7c74;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h261; din <= 32'hc0ef93e1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25e; din <= 32'h0956fd82;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20e; din <= 32'h356076aa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h233; din <= 32'h784f9af9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h001; din <= 32'h2fe133d4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h156; din <= 32'haaf759eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24d; din <= 32'hfa8dbf32;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h272; din <= 32'h5e104244;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h286; din <= 32'h782ed5f1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c2; din <= 32'he3a54c74;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3de; din <= 32'hb22a0fe2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b9; din <= 32'hd11dacdd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h276; din <= 32'h0c52db18;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18e; din <= 32'h3f971f19;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12d; din <= 32'h11724b1a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h118; din <= 32'h97583f86;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d4; din <= 32'h82ef8d83;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04e; din <= 32'h7a0efb8e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d9; din <= 32'had7f5b3d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h299; din <= 32'h93e39363;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h026; din <= 32'h53cb1df6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b4; din <= 32'ha4e6b621;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15b; din <= 32'h43aebccb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bd; din <= 32'hff8d7877;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h341; din <= 32'h5e35c2bf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ed; din <= 32'h02b3a2ad;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h367; din <= 32'hf31e250f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h063; din <= 32'hd9adc794;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09b; din <= 32'h7b2dea74;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ca; din <= 32'ha9ce2bf1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a4; din <= 32'h6fd627f7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33b; din <= 32'hd8e04bf4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h373; din <= 32'hb5741ee8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19b; din <= 32'hffeab59c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03f; din <= 32'h647f6803;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h114; din <= 32'hf033dfc2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h244; din <= 32'h8aeb5cbc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h351; din <= 32'h2339874a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06c; din <= 32'hbb9a2154;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cd; din <= 32'hf20fff71;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h267; din <= 32'hc57058a8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14b; din <= 32'hb3a9381e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h190; din <= 32'ha621b0e3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h254; din <= 32'h71443173;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h365; din <= 32'ha6dfc392;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2de; din <= 32'h68061317;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h047; din <= 32'hf45dd8aa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c6; din <= 32'h9cf9579c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h307; din <= 32'h9cd37efb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f3; din <= 32'h1857106f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17d; din <= 32'h8cffcae1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06f; din <= 32'ha359ccd1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d0; din <= 32'h5111640e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h344; din <= 32'h5fc57074;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h315; din <= 32'hf30552d2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h191; din <= 32'h7443e6b7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d5; din <= 32'he02a77d8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h302; din <= 32'h7cb01df0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c0; din <= 32'h920479b7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2af; din <= 32'h1a5667b9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ea; din <= 32'h118ab441;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f0; din <= 32'ha0d4eb91;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e2; din <= 32'h03620560;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e4; din <= 32'h7ce5caa2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e3; din <= 32'hb9139aed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ca; din <= 32'h2691f766;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h047; din <= 32'h5dd7f605;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3db; din <= 32'h44c4411b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a6; din <= 32'h54d1212f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ee; din <= 32'he43ce92c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h279; din <= 32'h19d4bb5a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3aa; din <= 32'h2fb585cc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h114; din <= 32'h7497fcd1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h076; din <= 32'h14db217c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h016; din <= 32'h0c36d507;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a5; din <= 32'hd11145fd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h101; din <= 32'h3ed6f611;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h068; din <= 32'h1e38d9be;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h089; din <= 32'h5b961ec6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39c; din <= 32'hc0ca3599;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d2; din <= 32'hffc92796;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01d; din <= 32'h74022867;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e0; din <= 32'haf76a2e8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h231; din <= 32'h77f71e45;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d0; din <= 32'h7fcf7779;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h259; din <= 32'h93c1a337;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29f; din <= 32'h62fdbee9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h045; din <= 32'h872f3420;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c9; din <= 32'h4badc6d9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d6; din <= 32'hf6c05d5c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16b; din <= 32'hcfae1995;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cb; din <= 32'he1e42201;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3de; din <= 32'h0d864da9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e3; din <= 32'ha8f59c85;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21e; din <= 32'h16e17dbe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h204; din <= 32'h8358b7c1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h181; din <= 32'hb10f2424;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e7; din <= 32'h11aa2665;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06b; din <= 32'h5bce322d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f1; din <= 32'h09d01d32;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30e; din <= 32'hb1269772;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h188; din <= 32'h04aa7adc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2fa; din <= 32'h854fbab7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f3; din <= 32'he0ba2ef4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h376; din <= 32'hec68bb08;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38d; din <= 32'h977342b1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c0; din <= 32'hf6da5874;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0df; din <= 32'h553d1827;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a6; din <= 32'hfcc9a2d2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h230; din <= 32'h923886dd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cd; din <= 32'h4ca734a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a2; din <= 32'hdf7c77da;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06f; din <= 32'h09a8efcb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h296; din <= 32'h3814ea4e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28e; din <= 32'h0a5aeaea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h076; din <= 32'ha761fe45;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b1; din <= 32'h78ffe4dd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22b; din <= 32'h56c456d3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h302; din <= 32'hfc418b41;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h241; din <= 32'h3f73b2cf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2fa; din <= 32'h50959516;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h000; din <= 32'hdb21b938;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h221; din <= 32'h4bc47691;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10a; din <= 32'h11210e12;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06d; din <= 32'h6adbd41a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01f; din <= 32'h3ad58e26;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h228; din <= 32'ha65f2cc9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ea; din <= 32'h75f6120e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h164; din <= 32'hf00484ee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37c; din <= 32'h5ed1cbb2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h386; din <= 32'hde17650f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h346; din <= 32'h9dac1cee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c4; din <= 32'h018bc751;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h290; din <= 32'ha9cd2199;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a8; din <= 32'he895b63a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39b; din <= 32'h263a9af8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c2; din <= 32'h0b62379e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h230; din <= 32'hdac9cdae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h302; din <= 32'hf9dc1385;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h185; din <= 32'h0a450480;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h164; din <= 32'hf63b65ff;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c1; din <= 32'h330ff24c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h280; din <= 32'h9fbc384b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c3; din <= 32'h846121ac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a9; din <= 32'h6c2d0439;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h216; din <= 32'hc1049c42;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12e; din <= 32'ha9c08967;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h135; din <= 32'h36469f52;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f3; din <= 32'h783d0869;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h106; din <= 32'h2eb04f38;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h333; din <= 32'hf63ce537;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c5; din <= 32'haec598c3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h242; din <= 32'ha575bb09;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h284; din <= 32'h02e93320;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c6; din <= 32'h65a59807;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38f; din <= 32'hca7611fb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h184; din <= 32'hc5c9301f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ae; din <= 32'hb1ddcdae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fb; din <= 32'h7006785d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h328; din <= 32'h82e2a7ed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h139; din <= 32'h39c41687;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2fb; din <= 32'h31acaa12;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a0; din <= 32'h0103b519;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h180; din <= 32'hcfd15551;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h272; din <= 32'hc31bb146;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h154; din <= 32'ha179f3e4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ca; din <= 32'h742e68e5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3dd; din <= 32'h45a7cfba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e1; din <= 32'hd02660d9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25e; din <= 32'h11a276c9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b0; din <= 32'h5565e9a9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a1; din <= 32'hff1072ec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d7; din <= 32'hbb961acf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h326; din <= 32'hd64cf808;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27d; din <= 32'h1de54ebf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h092; din <= 32'h84fa338b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h262; din <= 32'h984b9d52;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21c; din <= 32'h18093e38;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h255; din <= 32'h82ff635b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33e; din <= 32'h03474975;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h120; din <= 32'h5d0438f8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h355; din <= 32'h42395d03;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07d; din <= 32'hf6de3d1a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14b; din <= 32'h04f8da86;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fb; din <= 32'h1fca7492;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h096; din <= 32'hc47bc270;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30d; din <= 32'h5d2527ca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34a; din <= 32'ha228b5f6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h274; din <= 32'hbda01df3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1dc; din <= 32'h66d08210;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07a; din <= 32'h021ada18;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h254; din <= 32'hd24b9e94;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h043; din <= 32'h990bebc7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h194; din <= 32'h5d352b98;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b0; din <= 32'h450f685d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e0; din <= 32'h11a230a3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h282; din <= 32'hcce9df78;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h018; din <= 32'h4e03d974;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h137; din <= 32'ha540d5c3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h267; din <= 32'hdc096e25;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12d; din <= 32'hd03a9d9e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cc; din <= 32'h18b2eefb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h073; din <= 32'hf94b90c8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d8; din <= 32'h20ff0fe7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b2; din <= 32'h5629e6e8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ef; din <= 32'he4bf88c5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32c; din <= 32'h07780b8e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h185; din <= 32'h19a66332;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cd; din <= 32'hf9aef8e3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d6; din <= 32'h6db98b00;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h397; din <= 32'h37e21f76;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h318; din <= 32'h8e778499;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ec; din <= 32'ha0469d6c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h355; din <= 32'hfd92f833;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h240; din <= 32'ha578cc9e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19f; din <= 32'h5d7a7fb6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h019; din <= 32'h020855ce;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a0; din <= 32'h16e5e423;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h140; din <= 32'h75a9f75f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39b; din <= 32'hd4f5f990;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h261; din <= 32'hb4b844c7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h262; din <= 32'h6fe383dc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e1; din <= 32'h3706a138;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32d; din <= 32'h26084e12;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b2; din <= 32'h9b26f2cc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36e; din <= 32'hbf7235c6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f2; din <= 32'h72b69886;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34f; din <= 32'h7e46a964;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ab; din <= 32'he5938b1d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fc; din <= 32'hae5cb85d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ae; din <= 32'h0e373536;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d5; din <= 32'h4626180d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d8; din <= 32'hbe090751;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h397; din <= 32'hf7e28911;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ae; din <= 32'ha91e0900;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a4; din <= 32'h553b5ef2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h079; din <= 32'h0aa77b16;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cf; din <= 32'h94abc87c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h218; din <= 32'h19d7e07e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b0; din <= 32'h1eecbd6c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h052; din <= 32'hafbb6896;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h194; din <= 32'h60c0f8a2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27e; din <= 32'h126c544a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c7; din <= 32'h4c079a18;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ec; din <= 32'h71af855b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h348; din <= 32'h6b908e33;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fd; din <= 32'he4f16360;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h146; din <= 32'h3b09ec20;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d2; din <= 32'hd3c57771;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e8; din <= 32'h018420e8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h157; din <= 32'hdc6d45f6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h370; din <= 32'hc90fa496;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35d; din <= 32'h6e9ba6f2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h097; din <= 32'h0683d2a1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08f; din <= 32'h4f7b9b59;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b6; din <= 32'hc2dfb6ac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a0; din <= 32'h5087d990;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h193; din <= 32'h16ea9eac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06d; din <= 32'hebe1d135;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f1; din <= 32'h69ff49b0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a9; din <= 32'h6027a3c6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cb; din <= 32'hecf14790;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h055; din <= 32'h1af33218;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a6; din <= 32'h1c3a6328;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d5; din <= 32'hb96f4c48;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h067; din <= 32'hfadbdf1a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h343; din <= 32'h1d0d3ef8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ce; din <= 32'hd845c3ae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h176; din <= 32'habbb7b98;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h137; din <= 32'h03377129;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b8; din <= 32'h9a9d949b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a1; din <= 32'h1833f4af;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0dc; din <= 32'hf64cd43a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h018; din <= 32'h2ec7ce60;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h161; din <= 32'h7dd653da;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f7; din <= 32'hf08b00e1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fd; din <= 32'hb0bac104;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09b; din <= 32'hd05a007c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h002; din <= 32'h90de1f71;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h078; din <= 32'h583a5a1d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h378; din <= 32'h99ec4093;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h217; din <= 32'h6e5ecc53;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e3; din <= 32'hde59e1d1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31e; din <= 32'h63ed88f4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3dc; din <= 32'h855df8ee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28a; din <= 32'h70a09256;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24a; din <= 32'h0626cb15;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h398; din <= 32'h4149d405;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e7; din <= 32'hf00e17b9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17b; din <= 32'h5d7bbf2e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c5; din <= 32'h7b7bdcc7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h050; din <= 32'hc4cc3cae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ea; din <= 32'he9867dd2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h083; din <= 32'hcea37d64;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bf; din <= 32'h50d19487;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bb; din <= 32'h9a1d42ce;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h201; din <= 32'h228d324e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h141; din <= 32'h7507a20e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0db; din <= 32'hb4009a42;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h153; din <= 32'hd8e5d45a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h059; din <= 32'h49878d4e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h051; din <= 32'ha1788e72;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h171; din <= 32'he7bf601c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31e; din <= 32'h3669643d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h224; din <= 32'h2638aabe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c3; din <= 32'h099fde23;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h212; din <= 32'h7adc1ef5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0eb; din <= 32'h6ddfd086;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19e; din <= 32'ha86d450d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18b; din <= 32'hba6dcbce;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06c; din <= 32'h147716f9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b5; din <= 32'hd999f7aa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h354; din <= 32'hd5f8ecad;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b4; din <= 32'h94e882f8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e5; din <= 32'ha255cc39;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f3; din <= 32'h1ba672fa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a8; din <= 32'h0b89f4f2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h109; din <= 32'hb043f2ee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c3; din <= 32'h566f74f4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h186; din <= 32'h78d97d15;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h350; din <= 32'habaa33b4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cb; din <= 32'h98039a67;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29a; din <= 32'h4cea8db8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h256; din <= 32'h3ddabe9a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17a; din <= 32'h38d69d78;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c0; din <= 32'h02b42a02;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10d; din <= 32'h2097846e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a8; din <= 32'h2412155c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h004; din <= 32'he5d77822;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h049; din <= 32'h523b5b4a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13b; din <= 32'h9d2a9a40;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h145; din <= 32'ha1f5b9f7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d6; din <= 32'h4144db09;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h132; din <= 32'heb5c21b2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38d; din <= 32'hd45d608d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23a; din <= 32'h8db87b5c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h344; din <= 32'hb8c077ef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h038; din <= 32'hce271587;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h244; din <= 32'h68ee81e0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e1; din <= 32'h2e650f2b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ac; din <= 32'hd8ebeec6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c8; din <= 32'h609e761c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a5; din <= 32'h6013eec5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38f; din <= 32'h276701e1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h375; din <= 32'h635a5ffd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e6; din <= 32'h158d7c54;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c3; din <= 32'h8a0655d7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h233; din <= 32'h837ea593;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h037; din <= 32'h39cd2a40;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f1; din <= 32'hca1dcfda;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2aa; din <= 32'h0bf43f21;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10f; din <= 32'h5359e8d7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fa; din <= 32'h2f6e255c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1da; din <= 32'he5fe6180;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34c; din <= 32'h269aae0e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h057; din <= 32'hdc50a4be;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e3; din <= 32'ha140a7a5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h055; din <= 32'hd2c7d9b3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23d; din <= 32'he1e03588;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22e; din <= 32'hee6a9e40;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c5; din <= 32'h667b698d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h168; din <= 32'h0732f029;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b9; din <= 32'h012f6806;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f5; din <= 32'h5e2b8fb7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h392; din <= 32'h31793dc4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31a; din <= 32'haa80558f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ac; din <= 32'hd906cc90;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27e; din <= 32'h4324dc50;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h233; din <= 32'h955a714a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h108; din <= 32'h493c25c3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h281; din <= 32'hcf7b8a37;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h073; din <= 32'hd6060c7d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d0; din <= 32'h08e02471;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h336; din <= 32'h15c9d9fd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h199; din <= 32'hd911906f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h188; din <= 32'h46bc5821;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h166; din <= 32'h44e2921d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h047; din <= 32'h46d4559f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21b; din <= 32'h1fa34d28;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h212; din <= 32'he8cf8b41;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26d; din <= 32'h9f0c630b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a9; din <= 32'h915c5119;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h276; din <= 32'ha83d8014;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0eb; din <= 32'h45631af8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h117; din <= 32'h6f1b96e7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h393; din <= 32'h9ee138e0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1db; din <= 32'hf9effb99;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21e; din <= 32'h9083934b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28d; din <= 32'ha0204760;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12f; din <= 32'h944f00d6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f6; din <= 32'h70eba396;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h093; din <= 32'h5dddb899;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h096; din <= 32'he61286f8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h024; din <= 32'hcd1d914e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h154; din <= 32'h78cdd772;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h019; din <= 32'h1989ef1d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35d; din <= 32'h5f6468e5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26e; din <= 32'h5cebdabe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c7; din <= 32'hfc9ea327;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h053; din <= 32'haee4a41b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b3; din <= 32'h5466db83;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c2; din <= 32'h92d82097;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36b; din <= 32'hca402b79;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h186; din <= 32'h7c90a43e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a1; din <= 32'h6bdb302d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a1; din <= 32'hf1cb3c22;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h392; din <= 32'h106d481a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f7; din <= 32'h8ae24815;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h310; din <= 32'h993264bb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18e; din <= 32'hb076b9a7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f4; din <= 32'hf931863f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h127; din <= 32'hcff4ce66;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b8; din <= 32'hd340863d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ad; din <= 32'hba75d249;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h226; din <= 32'hdbc6d267;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h214; din <= 32'h7b9e7bb5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1aa; din <= 32'h671fabf8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h187; din <= 32'h8db58d17;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38a; din <= 32'h3a5a7a90;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23b; din <= 32'h8ed53daf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33e; din <= 32'hdab207e0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29e; din <= 32'haec8fb1d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e9; din <= 32'hd37b5952;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d7; din <= 32'h865465cb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07f; din <= 32'hd5c0e5ad;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d9; din <= 32'hd3c8ef0a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a2; din <= 32'h2d7fa05c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h048; din <= 32'h8f7d195f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34c; din <= 32'h1d213ab6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a8; din <= 32'hfe0e4244;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39a; din <= 32'h815f182b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h392; din <= 32'he8b622f3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25d; din <= 32'h71ff4e6b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f8; din <= 32'h6a48804a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15d; din <= 32'hf9a17dd5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1dd; din <= 32'hda88cc04;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ba; din <= 32'h16b3ae8c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h134; din <= 32'h013d6bd3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h215; din <= 32'h9b34a14d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27b; din <= 32'he01f64ae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h038; din <= 32'h0cba5c1c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ab; din <= 32'h685d542a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e9; din <= 32'h6cd3591a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39b; din <= 32'heb9c6e55;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f8; din <= 32'h2937c152;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c0; din <= 32'h9548d31f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h280; din <= 32'h44242660;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a4; din <= 32'hd0377f79;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d6; din <= 32'h277585a7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e3; din <= 32'hbd12290d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32b; din <= 32'h5bbe0d01;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27d; din <= 32'he74748ff;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h347; din <= 32'h02ccbd5f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h312; din <= 32'hce64278a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f4; din <= 32'h73e66ffc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28f; din <= 32'hdc9053c0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h231; din <= 32'he3d7fce8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h208; din <= 32'h2e919026;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d2; din <= 32'h87beae82;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ed; din <= 32'hb70ff8fd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h361; din <= 32'h465dc868;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c5; din <= 32'h7f7cf733;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ed; din <= 32'hd4cef6b1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05c; din <= 32'h479d8639;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h396; din <= 32'hc40d0e5a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h110; din <= 32'h822a37e0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ce; din <= 32'he5721558;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24a; din <= 32'h72f155b9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0eb; din <= 32'hf87bafb2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c5; din <= 32'h60d28d37;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h213; din <= 32'ha9980d84;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ba; din <= 32'h071e4179;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h092; din <= 32'h3f2e1f7f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h308; din <= 32'h9b08c7db;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e0; din <= 32'h9ce79eaa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12b; din <= 32'h1c218f7d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f1; din <= 32'h91510d24;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a1; din <= 32'h731ea0ae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e8; din <= 32'hce4d1fae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13a; din <= 32'h274d4182;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11f; din <= 32'hd9009725;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14a; din <= 32'he2bd4537;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h020; din <= 32'h102fd8f1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h274; din <= 32'h8559e20c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h277; din <= 32'h2469a21f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h086; din <= 32'h18f3d658;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a9; din <= 32'h35cae39e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ec; din <= 32'hd3f8d119;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b5; din <= 32'h5862c594;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06e; din <= 32'h3bc54b14;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25f; din <= 32'h13855603;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37c; din <= 32'h4d0e5777;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h326; din <= 32'he40ab879;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ed; din <= 32'hfb47f66c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06c; din <= 32'hec1427ab;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h114; din <= 32'he792883c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b4; din <= 32'h197b0e00;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h309; din <= 32'hc8a607de;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03e; din <= 32'h525a5b5a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b3; din <= 32'h703140a1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a2; din <= 32'h58303e6c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h142; din <= 32'hba846b92;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d4; din <= 32'h17f73e1b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30a; din <= 32'hc5ab64fe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15e; din <= 32'hc8030e6e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c7; din <= 32'h51f76923;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c1; din <= 32'hc21ac646;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bd; din <= 32'h62dc4757;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ce; din <= 32'hdc3cbe01;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h120; din <= 32'h851e6500;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ca; din <= 32'h805ace2b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07d; din <= 32'h599b91a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a1; din <= 32'hb8bec9e6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ae; din <= 32'he9e7c305;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b6; din <= 32'h70ac9452;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h389; din <= 32'h6019517f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3de; din <= 32'he66f00a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h341; din <= 32'h5895a1ef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h330; din <= 32'h03e306eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35f; din <= 32'hacf39607;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e5; din <= 32'hdc0a9e9f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e7; din <= 32'hb283d1fc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h081; din <= 32'hb782565d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03e; din <= 32'h8937f276;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cb; din <= 32'hddd1fe88;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c4; din <= 32'h869f93ea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h009; din <= 32'hddb9487a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d5; din <= 32'h2f4ff433;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31e; din <= 32'h45dccad3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09c; din <= 32'hffe2b3f3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3aa; din <= 32'h00b42eb9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14c; din <= 32'h1aaa4b3d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16b; din <= 32'h26a047f2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h290; din <= 32'h15676291;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02b; din <= 32'h42b938a9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f8; din <= 32'hbccd172c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h389; din <= 32'h6a0ef6cc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h184; din <= 32'h783b9f80;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09f; din <= 32'h6dce789f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03c; din <= 32'h598fda98;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25c; din <= 32'hc50b9c3f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12f; din <= 32'h8e30c8b8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06a; din <= 32'h592c1cd2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a9; din <= 32'hbc862da1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02c; din <= 32'h440b082c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3aa; din <= 32'h39aef79e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e8; din <= 32'h37b7b68d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h394; din <= 32'hffd03ee1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h194; din <= 32'h8f79bc1c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h116; din <= 32'h1bdcce30;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h148; din <= 32'h414e0fbf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f6; din <= 32'hdd60feeb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09a; din <= 32'h87104abf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0af; din <= 32'h5c8910f2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e8; din <= 32'hb4e67683;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36f; din <= 32'h97a37bbc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30d; din <= 32'hcb01be72;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f6; din <= 32'h3d42a23a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h098; din <= 32'h74d0d0e8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f7; din <= 32'hd406985f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01b; din <= 32'h22a8d198;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f8; din <= 32'he167d0b0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cd; din <= 32'h0f0bc7ad;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h169; din <= 32'he396e537;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h237; din <= 32'h1bcc12c4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e3; din <= 32'h45f5a2dc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h299; din <= 32'h17ef9b1f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h066; din <= 32'h998aec39;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h288; din <= 32'h085c5b7e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h117; din <= 32'hecc76ad4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b3; din <= 32'h846f9e13;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24a; din <= 32'h322de95f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d6; din <= 32'h76c6ff30;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19b; din <= 32'hf41ccc73;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ce; din <= 32'h44ea7650;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cc; din <= 32'h42a22265;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29a; din <= 32'ha2bebbef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fd; din <= 32'hf13910dc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h155; din <= 32'h015e6bf9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cd; din <= 32'hb44050c6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23d; din <= 32'h6c760d04;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f2; din <= 32'hce1f148b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24a; din <= 32'hbaf92b36;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h117; din <= 32'h263a2ddd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b4; din <= 32'h3ca09808;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21e; din <= 32'hd4802789;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ed; din <= 32'hc52cafb4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f9; din <= 32'ha246a070;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c3; din <= 32'h3835a841;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03b; din <= 32'h5ceb2ec9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38b; din <= 32'hbc5d3dcf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ce; din <= 32'h6ced761f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h088; din <= 32'ha0612c92;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h040; din <= 32'h2f8dcb56;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h212; din <= 32'he88be3a7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b2; din <= 32'hd8d54316;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26a; din <= 32'h49e7a1ab;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h113; din <= 32'h376a6abb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h275; din <= 32'h2f4ed3b7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cd; din <= 32'h06afd82b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h120; din <= 32'hf425a25a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21d; din <= 32'h1a714e90;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31d; din <= 32'hc7ab1676;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h063; din <= 32'h803c1722;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bb; din <= 32'he10f1dc2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h177; din <= 32'h2f85f92f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h281; din <= 32'hade96823;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h386; din <= 32'h9573eceb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h150; din <= 32'h2c4717bb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d1; din <= 32'he4fafe4e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37e; din <= 32'h841b73b7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h397; din <= 32'hcf0f8671;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d3; din <= 32'h68b6a52f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1dd; din <= 32'h57fef2fa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13a; din <= 32'h566645a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24d; din <= 32'h13b243dc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h235; din <= 32'had3ed8b9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15c; din <= 32'h865d9faf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29d; din <= 32'h20dfd7f7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e3; din <= 32'hb107d14e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f6; din <= 32'h0e18276f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09f; din <= 32'ha8195c7b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h020; din <= 32'haecedfa0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h342; din <= 32'h90cddf0e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b2; din <= 32'h9e8345ca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e3; din <= 32'hf21016c5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h320; din <= 32'h0e8f8e7c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h228; din <= 32'hd35da938;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01e; din <= 32'h17eebf07;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h211; din <= 32'hc01e450f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b1; din <= 32'hc1deb3bb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37d; din <= 32'h9359e4f5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03f; din <= 32'h2afcacc7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h064; din <= 32'h28ab8fd1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h311; din <= 32'hef89b964;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ec; din <= 32'h55ed66f0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h396; din <= 32'h601e9884;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26c; din <= 32'h22841247;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h370; din <= 32'h62bca218;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h060; din <= 32'hbb3e3eb3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e0; din <= 32'h824b27b0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ce; din <= 32'h8306c4fb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28c; din <= 32'h50d909fe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h107; din <= 32'hcb88d7f7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h145; din <= 32'hd98a576a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1df; din <= 32'h9db42f14;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f1; din <= 32'h649d081a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c2; din <= 32'hb170e537;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bc; din <= 32'he0734877;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h387; din <= 32'ha8834337;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h017; din <= 32'hbff9d0fd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b4; din <= 32'h223e2fa5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d7; din <= 32'hf70d6980;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h379; din <= 32'h3aa90b4a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32a; din <= 32'hf8bc2bae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h196; din <= 32'h29f25f67;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a8; din <= 32'h8076907f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25c; din <= 32'hc99ba74f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c7; din <= 32'h7dd6c7c9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h213; din <= 32'h685fb476;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c9; din <= 32'hf37744b4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h077; din <= 32'h5a7908f6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h309; din <= 32'h887b20c1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h057; din <= 32'h72b54bbc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b7; din <= 32'hb4e10d95;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h265; din <= 32'h0a63ca36;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h025; din <= 32'h0523e690;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h210; din <= 32'he4b2700b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e1; din <= 32'h6c6a3c41;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ea; din <= 32'h88dcd66f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h082; din <= 32'h696fc711;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e1; din <= 32'hfc6f5c16;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19c; din <= 32'h65372fa4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00c; din <= 32'hc649e7a8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37d; din <= 32'h8b42da79;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b1; din <= 32'hd4a7c9ab;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h058; din <= 32'hc1e8f0f4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h212; din <= 32'hdfc800af;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h221; din <= 32'h63875884;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h290; din <= 32'hf4e4e1bc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ca; din <= 32'h74356675;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h248; din <= 32'h61ebf82e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h398; din <= 32'h661bda5d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13f; din <= 32'h169863e6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00c; din <= 32'h033fa984;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h036; din <= 32'h98a7a4de;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fc; din <= 32'hf54d8312;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h016; din <= 32'h91ee8daf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2aa; din <= 32'h37b1cdf8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h067; din <= 32'h85cffd70;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h326; din <= 32'h387def76;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f1; din <= 32'h3f7f4208;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h267; din <= 32'hdc0944f4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ef; din <= 32'h31993133;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a9; din <= 32'hc7f3af1f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29a; din <= 32'he4541026;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h024; din <= 32'h15022e93;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f8; din <= 32'hcfe68698;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33e; din <= 32'hfa34cb2b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bb; din <= 32'h30631deb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d9; din <= 32'h9418e453;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05b; din <= 32'he546b508;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d8; din <= 32'hb225d53a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f2; din <= 32'hfc840ce8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ca; din <= 32'h522415cd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13b; din <= 32'h2f1bd442;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26c; din <= 32'hcde8ab42;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b4; din <= 32'h57e692df;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h278; din <= 32'h4b9486be;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h394; din <= 32'h022d056e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h155; din <= 32'h1281d494;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h334; din <= 32'hf3d0c0de;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h165; din <= 32'hdf4bd731;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16e; din <= 32'hd5de5e1f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h170; din <= 32'hcbc634b7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h205; din <= 32'h55bf05fa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a8; din <= 32'h0027fbe5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h171; din <= 32'hc4de7e6d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h215; din <= 32'h5a0823db;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27e; din <= 32'h8083a629;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ea; din <= 32'hef948670;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d5; din <= 32'h513bfe32;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34b; din <= 32'h3a856071;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ac; din <= 32'h19d67075;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h178; din <= 32'he4f978ce;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e7; din <= 32'h492c062e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c5; din <= 32'h0fcc38e0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h343; din <= 32'h5ea80c82;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2da; din <= 32'h47960fef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f5; din <= 32'h494d253a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h335; din <= 32'h999f2251;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e4; din <= 32'hd8337f3d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f5; din <= 32'h823bc748;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h356; din <= 32'h4102ddaf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c9; din <= 32'h1130cbad;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08a; din <= 32'h87ba1d74;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c5; din <= 32'h7dbeac49;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24d; din <= 32'h744abfa6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h198; din <= 32'hbf3d5fe3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d0; din <= 32'hec4b9b2f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h032; din <= 32'h4e14fe16;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ac; din <= 32'h5eda0bf0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h220; din <= 32'h2c751a38;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h107; din <= 32'heca6086e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cd; din <= 32'hdc6a8df7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b6; din <= 32'he2d4dd7e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h172; din <= 32'h0b2dda2f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h063; din <= 32'h0e576098;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3df; din <= 32'h8bde95ec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35c; din <= 32'hd86920fc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28b; din <= 32'h4f4f8132;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h203; din <= 32'h036797f9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19f; din <= 32'he780a24f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02e; din <= 32'h17472b32;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09e; din <= 32'h10f1d9d7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h090; din <= 32'hbabd844d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02f; din <= 32'hdafa231b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h340; din <= 32'heccd1b25;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c0; din <= 32'hb8cd985e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ef; din <= 32'h00e4f8c1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12a; din <= 32'h0009123d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b5; din <= 32'h408c62e2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ce; din <= 32'h4d7f4e7f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13c; din <= 32'he463c715;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h355; din <= 32'h788a871f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h050; din <= 32'h42788f57;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e3; din <= 32'h80e4269f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25f; din <= 32'h13ba4fe8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24f; din <= 32'h1bf537c7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23c; din <= 32'hc86d0516;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h211; din <= 32'h1ade55b0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2fd; din <= 32'hdde4a830;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f7; din <= 32'h45dcd29e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24f; din <= 32'h4f859f2c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d4; din <= 32'h3e9ab902;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05a; din <= 32'h09697523;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h324; din <= 32'hddaf015c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31c; din <= 32'h7271a325;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d1; din <= 32'h5d8c065f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h328; din <= 32'hbc34b59f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f4; din <= 32'hab3fd5a9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h326; din <= 32'h18ebffac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h098; din <= 32'h948f9920;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c5; din <= 32'hf9817182;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h302; din <= 32'he2007b3d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25c; din <= 32'hb5a1de69;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f1; din <= 32'hbfe76a65;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h052; din <= 32'h18bfc684;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d4; din <= 32'h65d594d0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d7; din <= 32'h303f7b9b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f8; din <= 32'hf24933ae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24b; din <= 32'h2e7dbf84;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09c; din <= 32'h1c13e40b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ed; din <= 32'h3a9ef49b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h386; din <= 32'h712fb946;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09a; din <= 32'h85fb19dc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12f; din <= 32'hc0ba2963;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cf; din <= 32'h1c7faeb7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39a; din <= 32'h08017ee4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08b; din <= 32'h76daad98;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cd; din <= 32'hfbd9cdea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h082; din <= 32'haea0798f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b2; din <= 32'h518547cb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39c; din <= 32'hf944778b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01d; din <= 32'ha7f161e3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h061; din <= 32'h83d14294;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2fa; din <= 32'hfbf9897c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h061; din <= 32'h9566e138;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d6; din <= 32'h0b5eaf9f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a6; din <= 32'he41e0ff6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h017; din <= 32'h859d057b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bb; din <= 32'h2b60c07a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08a; din <= 32'hc49a949f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20f; din <= 32'hb632480d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h329; din <= 32'heb69bc63;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cb; din <= 32'h3b0f0b78;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ec; din <= 32'h0759c0db;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ae; din <= 32'h5b57a3a5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h072; din <= 32'h40f201a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a5; din <= 32'h72015edd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b8; din <= 32'he7c27c6f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06a; din <= 32'h94404db5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h324; din <= 32'h0b567cc1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d0; din <= 32'hc15fd8a5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3df; din <= 32'h9139b3e2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d4; din <= 32'hd75f471a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d1; din <= 32'h4a61972b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h014; din <= 32'h27e249df;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a3; din <= 32'hdc11dc74;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h245; din <= 32'h997ddf32;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3aa; din <= 32'h4c4bf4eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h370; din <= 32'h5fd3db0c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e4; din <= 32'h80ac07ea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h377; din <= 32'hcc6a6a81;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3eb; din <= 32'h5d25cbc9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bf; din <= 32'h25a9862e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19c; din <= 32'h64401ea7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24d; din <= 32'h14d77138;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22c; din <= 32'h496c4e6f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e9; din <= 32'hd42d74c3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h300; din <= 32'h893a6248;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c5; din <= 32'h967b416c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a7; din <= 32'h2da85ea7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e6; din <= 32'ha451901f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1be; din <= 32'h993a1ee8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h275; din <= 32'h0ccf7264;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b5; din <= 32'hab09c430;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ad; din <= 32'h9b8d8409;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h013; din <= 32'hd94d3e26;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h204; din <= 32'h016fccbc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h162; din <= 32'h3ec582e4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ab; din <= 32'h367ce792;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h260; din <= 32'hf8a705ed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3da; din <= 32'hd1b358a4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h005; din <= 32'h3c617a84;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b3; din <= 32'h38cdb78a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h222; din <= 32'h2ff80a37;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h259; din <= 32'hfe3cae0b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h028; din <= 32'h5ed91267;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h136; din <= 32'h8114624b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bf; din <= 32'h7adf5de7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h034; din <= 32'h7eae1337;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h192; din <= 32'hdfb92bfa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h137; din <= 32'h344c2f7d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2af; din <= 32'hbf48e9fc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ee; din <= 32'h2c06f92b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01d; din <= 32'hd5021dcf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07a; din <= 32'h50c3b0c4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e1; din <= 32'h67a0bf7f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d6; din <= 32'had4e321c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h165; din <= 32'h09e1fff8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38d; din <= 32'h2a01d04a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d2; din <= 32'hfa728407;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h170; din <= 32'hb10ae91b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h396; din <= 32'h7de7a496;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06a; din <= 32'hf5682e12;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h001; din <= 32'h26ffa924;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fe; din <= 32'h42232db5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h046; din <= 32'h6abe4ad5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e9; din <= 32'h135dda5b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2da; din <= 32'h67121c45;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25f; din <= 32'hf717d8cc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f8; din <= 32'h36ab80d9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34a; din <= 32'h810ecb88;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f3; din <= 32'h879c9ec0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f4; din <= 32'hb4c4f2b5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h073; din <= 32'h9f795c24;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d1; din <= 32'h7adf99d5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29a; din <= 32'h352e8aad;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a3; din <= 32'h9f5f482a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h030; din <= 32'h751864e0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a8; din <= 32'ha0a4f984;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h380; din <= 32'h59fbfdd8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a3; din <= 32'hc532c5a7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d9; din <= 32'h394a0992;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17b; din <= 32'hfe1006b9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28c; din <= 32'h0372ea0c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h244; din <= 32'h209af7de;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c2; din <= 32'h28265ecd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h114; din <= 32'h6ba16671;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f7; din <= 32'hb34b1c27;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h027; din <= 32'he87ca226;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0be; din <= 32'hb9098c5a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h085; din <= 32'hc791bc0e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27b; din <= 32'h8127b755;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32b; din <= 32'h5dc98d01;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h253; din <= 32'h54b5f9c4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e9; din <= 32'h037cc291;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f8; din <= 32'hc2cfdaf3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0da; din <= 32'hca107ca1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h043; din <= 32'h2467f6b6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34d; din <= 32'h2d958adf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d7; din <= 32'h09b64d3b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h257; din <= 32'h97631443;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h397; din <= 32'h210827f5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0df; din <= 32'hae265df2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33f; din <= 32'h617088eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23c; din <= 32'h56ff9077;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19a; din <= 32'h6d67b877;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h179; din <= 32'h172132e2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ef; din <= 32'hf764c8ca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h196; din <= 32'h08b0ec7c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f0; din <= 32'h84cdc259;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20c; din <= 32'h64284b08;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b2; din <= 32'h979b385b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b9; din <= 32'h855e2c49;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h125; din <= 32'h0aa5f38f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c9; din <= 32'h3777a269;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3db; din <= 32'h170022de;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21b; din <= 32'he6a84f46;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18b; din <= 32'h1bb7c224;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h007; din <= 32'hc4f10f5a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h378; din <= 32'hd21f35e7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37b; din <= 32'h7adcd543;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h018; din <= 32'h51b7074b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e8; din <= 32'h62da4841;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07d; din <= 32'h59663ec1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08b; din <= 32'hbf0745b8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16b; din <= 32'h68b27a2d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h217; din <= 32'h538fba62;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34f; din <= 32'h99507cbb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h212; din <= 32'h669bd5d2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h266; din <= 32'h7562be1d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h120; din <= 32'hdafc01f1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cd; din <= 32'h51bb65e0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h374; din <= 32'h0c407d63;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h054; din <= 32'hfa3b2f81;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bf; din <= 32'ha374b872;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h336; din <= 32'h340b9c54;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h398; din <= 32'h93e22b25;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h247; din <= 32'h777ce39c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h285; din <= 32'hb12a31ab;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f6; din <= 32'h761d911d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h275; din <= 32'ha6f7186c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24f; din <= 32'h52acf574;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h345; din <= 32'h553fee7d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h038; din <= 32'h2e1e35f1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ef; din <= 32'h169916a9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e7; din <= 32'h5d60f0a8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1db; din <= 32'h879e4245;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h169; din <= 32'hc8a58226;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d1; din <= 32'h1ba771cb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b7; din <= 32'hafd6d69d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b7; din <= 32'h99d10771;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f9; din <= 32'h0561bfb7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ae; din <= 32'h79368e2d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h354; din <= 32'h558e1fb8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c8; din <= 32'h4f5e6b05;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h038; din <= 32'hf9f372f9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11e; din <= 32'hca80acce;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f1; din <= 32'h29f0fce5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ec; din <= 32'h452d6c09;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01a; din <= 32'h1f91758d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33c; din <= 32'he1b4e294;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h103; din <= 32'hf80b867c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ce; din <= 32'hbcbbe715;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h371; din <= 32'h13ba8829;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h343; din <= 32'h599de3c5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24f; din <= 32'haa3cac4d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h326; din <= 32'h7b6c98a8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08c; din <= 32'h60aef431;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a2; din <= 32'h000194e5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h347; din <= 32'h903ee439;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f8; din <= 32'h1884eabc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h283; din <= 32'h33381d2e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h097; din <= 32'h40eed09b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h148; din <= 32'hf3b26b24;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d0; din <= 32'h86ef6ba9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e4; din <= 32'h3c6fd5e2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05c; din <= 32'h68f00f10;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04a; din <= 32'h9b2478f2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h347; din <= 32'h6cf346ed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h257; din <= 32'hae4c7293;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18e; din <= 32'ha21e6a10;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36d; din <= 32'h20105d2d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19e; din <= 32'hac970942;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b0; din <= 32'h83ac9018;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h264; din <= 32'h4bedd6de;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h344; din <= 32'hd26593fb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h336; din <= 32'h5ada8c6a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d6; din <= 32'h8f285c0c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17f; din <= 32'h694001aa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h070; din <= 32'ha8ac5894;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h241; din <= 32'hbaf43db4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h297; din <= 32'h8871bdce;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16f; din <= 32'hd0ef2de9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h243; din <= 32'h2b96dcb2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h141; din <= 32'hb0699e1b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c1; din <= 32'h02c49109;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h042; din <= 32'h4e0ea64b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c3; din <= 32'h2c960325;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h002; din <= 32'h3d37b78e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39a; din <= 32'ha1b026ac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h369; din <= 32'h1856cf63;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h165; din <= 32'hde91d0b9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1dc; din <= 32'hd7e374c8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h110; din <= 32'h71726568;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f2; din <= 32'he93be9ee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h352; din <= 32'hbfb2c3ed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cc; din <= 32'he5b34f25;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h323; din <= 32'h160daa80;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34d; din <= 32'h20c446ce;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19c; din <= 32'h6b676f97;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e1; din <= 32'hc326e951;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h090; din <= 32'h5c758224;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h238; din <= 32'h8a49a1bc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h061; din <= 32'h2fad9247;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d3; din <= 32'h7d207215;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ad; din <= 32'ha2171ab9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h162; din <= 32'hb7d71654;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33a; din <= 32'hf471558f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h041; din <= 32'h389a286b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28f; din <= 32'h874e6cee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h114; din <= 32'h516285b4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39b; din <= 32'h43debcf5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c7; din <= 32'hc14ab2e3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c4; din <= 32'h3a2964bc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d7; din <= 32'ha383530b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c3; din <= 32'h72c02aea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07d; din <= 32'heca71a07;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a3; din <= 32'hfb616584;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c6; din <= 32'hd0e6feeb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2fa; din <= 32'hea1a1875;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f7; din <= 32'h86d820ee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h257; din <= 32'h95575fac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h208; din <= 32'hadf2eff2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h136; din <= 32'h0c310eea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c3; din <= 32'he3b8d009;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a7; din <= 32'h83bfa862;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e6; din <= 32'heb403a4a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h285; din <= 32'he6b31a2b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08c; din <= 32'hd9acdb7b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e7; din <= 32'hcbfe7fb6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c4; din <= 32'h7bc8057b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34c; din <= 32'haf2cea8b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ea; din <= 32'ha4f29f00;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h341; din <= 32'h5da37e61;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h334; din <= 32'h41d31759;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h348; din <= 32'h7c0bdb7e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0af; din <= 32'h70f346c8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19b; din <= 32'h95d16941;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c8; din <= 32'he7271a16;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h021; din <= 32'h7c87924e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1aa; din <= 32'h6c3881b5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bf; din <= 32'h2effeeba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h221; din <= 32'h12c54f40;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h218; din <= 32'h6c61b096;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25f; din <= 32'haa48a299;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b5; din <= 32'h5fa4b0cf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10b; din <= 32'h6dee7b1a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h064; din <= 32'hde015cd2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17d; din <= 32'h75848269;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h319; din <= 32'h01e61e4e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19c; din <= 32'h2b5a2544;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cd; din <= 32'h7edb95d8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h125; din <= 32'h2b328231;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23e; din <= 32'hf856ff14;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fe; din <= 32'h60cb95a9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15e; din <= 32'ha048d064;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f5; din <= 32'h8df9f914;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c9; din <= 32'h8ca59d29;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h018; din <= 32'h3ca09f1d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06e; din <= 32'he2f418df;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h031; din <= 32'ha172f6c5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2db; din <= 32'h41c1ef3f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h149; din <= 32'h47815987;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bf; din <= 32'h28255ed1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06b; din <= 32'h46ef2bd9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h340; din <= 32'h66ac8452;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h279; din <= 32'h89ec1388;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36f; din <= 32'h96d5ae2e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h025; din <= 32'ha9f86644;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16e; din <= 32'h91ae7c88;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f5; din <= 32'h344186e1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33e; din <= 32'hda730182;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h303; din <= 32'h0bff13b0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00c; din <= 32'h54a6447d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37e; din <= 32'h2bfa749a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h090; din <= 32'h4d94e1b4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h307; din <= 32'h74e12f0a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h394; din <= 32'h6318a868;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ae; din <= 32'hea5351d0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h179; din <= 32'h5a471c30;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d6; din <= 32'h92af27ea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e6; din <= 32'h7bb6bb6b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h287; din <= 32'h256e7770;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h242; din <= 32'he1a7592d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h303; din <= 32'hab0fe992;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h389; din <= 32'h3b7a11a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1dc; din <= 32'h554eadf0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ce; din <= 32'h989f37ef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ef; din <= 32'hc7f4d657;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ea; din <= 32'h147611f9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d7; din <= 32'ha5cc485d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a6; din <= 32'h57f7aa4a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b9; din <= 32'h30180c66;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04d; din <= 32'h19b23327;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39a; din <= 32'hae8f3368;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d9; din <= 32'he84e978f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f8; din <= 32'h8031123d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e7; din <= 32'h02cbffa0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a6; din <= 32'h8f26d4cd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h373; din <= 32'hfe1db039;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cc; din <= 32'h8eabc67d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3dd; din <= 32'h4702ebfd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31c; din <= 32'h3784a79c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33e; din <= 32'h1bc7ebb9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h357; din <= 32'h6fa3e156;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ac; din <= 32'h268c0575;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33e; din <= 32'h74810b41;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20f; din <= 32'h550e11a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c5; din <= 32'h1ff903d7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11b; din <= 32'h09369cb1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h114; din <= 32'hfbdaff10;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h183; din <= 32'h04348224;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h140; din <= 32'h673643bf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0dc; din <= 32'h191dc099;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11f; din <= 32'h7c44539e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06a; din <= 32'ha147f332;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b3; din <= 32'he20ddaf6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h056; din <= 32'ha31c1236;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h039; din <= 32'h4ed04b02;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h290; din <= 32'hd9ea33e0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h283; din <= 32'h5067476b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03b; din <= 32'h5df56d90;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h015; din <= 32'h06f84b89;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e1; din <= 32'hbbc8e17c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h306; din <= 32'h2487bf95;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c2; din <= 32'h7d43e286;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ea; din <= 32'ha6e6a8ea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bf; din <= 32'h630dfd68;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16d; din <= 32'h5d30e9d2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h241; din <= 32'h2df6d895;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e1; din <= 32'h93e63b24;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b3; din <= 32'ha321f45f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a1; din <= 32'h3d49b2a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h266; din <= 32'h0d94f903;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h153; din <= 32'h86b3fd03;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12e; din <= 32'hfec6f3ba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h316; din <= 32'hd9aabee0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e0; din <= 32'h7fe51109;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h080; din <= 32'h4520f9af;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f9; din <= 32'h3040187c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34b; din <= 32'he19bad28;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h220; din <= 32'ha99a3571;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h206; din <= 32'hbc1ea937;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h173; din <= 32'hddbe3ebf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h356; din <= 32'haf1a7402;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f3; din <= 32'hc7d76f3d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38c; din <= 32'h5e166160;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h314; din <= 32'h4ae2eb97;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1de; din <= 32'hc440d647;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h393; din <= 32'hb3e7dbf9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h242; din <= 32'hb88c8ad5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h210; din <= 32'h019066d2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h304; din <= 32'hb4042eb1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34f; din <= 32'h8105ac67;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fe; din <= 32'h55af1473;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2fc; din <= 32'ha5bfe8c0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b3; din <= 32'had1f69d8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ff; din <= 32'heb5d52af;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h136; din <= 32'hf98ab63c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a2; din <= 32'h7ed0fa92;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h116; din <= 32'h48a9f377;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h285; din <= 32'h1fa15806;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h227; din <= 32'h019b24b1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12d; din <= 32'hc689e4bd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fc; din <= 32'h7e786a08;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ad; din <= 32'h1cf7f80d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h265; din <= 32'hd23f149a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h365; din <= 32'hefceae8f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f4; din <= 32'h68927f0d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h357; din <= 32'hda31bc6e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ab; din <= 32'hb74ef796;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20e; din <= 32'h2864974a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c3; din <= 32'hc9dff106;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h244; din <= 32'hd380f64b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h169; din <= 32'hb291f1ba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h092; din <= 32'h0e5087e7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h233; din <= 32'hadd47ff7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e8; din <= 32'hbc48b25e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19a; din <= 32'ha4bc309d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d4; din <= 32'h7b541b52;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35a; din <= 32'hdc1bf089;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h105; din <= 32'hc7f12b8c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12e; din <= 32'ha0775196;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e3; din <= 32'h91b17000;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h354; din <= 32'hf9dd98d7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c6; din <= 32'hc3458a76;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h318; din <= 32'h32d8ba19;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h144; din <= 32'h4a0a7867;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h215; din <= 32'h1e3d32c3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h117; din <= 32'h16b51c1a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h151; din <= 32'h24f8f496;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29c; din <= 32'hd2919c65;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f8; din <= 32'h1f1fb1bd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b7; din <= 32'he3d5bb4d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h109; din <= 32'h79ef0a01;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ec; din <= 32'h4461623c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3eb; din <= 32'hd3f9df57;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h313; din <= 32'h7a563224;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h372; din <= 32'h391db616;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h066; din <= 32'h403c56f9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07b; din <= 32'h58ea92d1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h394; din <= 32'h18e324b2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19c; din <= 32'h0288bb39;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3de; din <= 32'hc36c3a0c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a2; din <= 32'h2c40a4e3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f6; din <= 32'h7a1e6312;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h293; din <= 32'h7e1f3e30;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18b; din <= 32'hd28d4b45;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h338; din <= 32'hf9c480a8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ad; din <= 32'h84c74d77;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18d; din <= 32'h6407f718;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ab; din <= 32'ha51edfdf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h168; din <= 32'hdf17bb17;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f5; din <= 32'h183765b3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22f; din <= 32'hf18156f4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h094; din <= 32'hff378945;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h096; din <= 32'hc6edad8b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h090; din <= 32'h9c04c230;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cb; din <= 32'h04e7fda8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h219; din <= 32'he7433f9e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02d; din <= 32'h56b8256d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06f; din <= 32'h1566531d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f2; din <= 32'h6a49dbf3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h347; din <= 32'h42700ef4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13b; din <= 32'heb4ce886;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h293; din <= 32'h20732552;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1da; din <= 32'hbd899a38;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h184; din <= 32'hd63ece50;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05c; din <= 32'h46bce4b9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c2; din <= 32'ha5b40177;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19d; din <= 32'h0e388e2a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h063; din <= 32'h713e1ec9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h323; din <= 32'hd7424bd7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h203; din <= 32'hc49dd47d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21c; din <= 32'h4c5db713;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h105; din <= 32'h6e41ffc9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22d; din <= 32'h46468efc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h228; din <= 32'h4a8f59ab;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03b; din <= 32'hfa986720;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h309; din <= 32'h14ba8957;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ac; din <= 32'h822e2065;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h315; din <= 32'hff0af541;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h014; din <= 32'hfa4d1a98;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b0; din <= 32'h6909c9cc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a6; din <= 32'hf2ae557f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a2; din <= 32'h704152f0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e0; din <= 32'hfa0e5cb9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h116; din <= 32'h1185fa74;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31b; din <= 32'h7a7b6ad3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h245; din <= 32'h55f25bbb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h235; din <= 32'hc06d95f0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h217; din <= 32'h6dbcf955;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b3; din <= 32'had995315;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11e; din <= 32'h8829b80f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14b; din <= 32'h8e91cecc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h101; din <= 32'hc6559227;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h381; din <= 32'h90a25cf9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h232; din <= 32'h8327f5e4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h313; din <= 32'h0a24a803;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h056; din <= 32'ha5386420;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3be; din <= 32'h78778a4d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29a; din <= 32'h7aabd178;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h221; din <= 32'h6eca5fbf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h044; din <= 32'h85b0d98a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a2; din <= 32'hbd99974b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a5; din <= 32'h1cf2af65;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f2; din <= 32'h2b11d821;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04c; din <= 32'h5cd2052f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h358; din <= 32'h22e3dcd9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b1; din <= 32'ha81038fc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h226; din <= 32'hb60f4728;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39d; din <= 32'h7be6e06d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27a; din <= 32'hd453d4d5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d2; din <= 32'h348c84cc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h287; din <= 32'hf1e245f1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f4; din <= 32'h5004c0e2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c4; din <= 32'h60f48b9c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h070; din <= 32'ha6c70842;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20d; din <= 32'h6ceaec7c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ce; din <= 32'h4680c7e4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07a; din <= 32'h0c98025c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00a; din <= 32'h82979e5d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e2; din <= 32'hf68c4329;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h022; din <= 32'h8ab0d844;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12d; din <= 32'h0af8ed30;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bf; din <= 32'h0de67d4f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h157; din <= 32'h654c79c2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h174; din <= 32'hbc062e76;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h079; din <= 32'h42009b85;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b8; din <= 32'he66466bc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3af; din <= 32'he780ff9d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04b; din <= 32'hba740356;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2af; din <= 32'h0a590414;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a1; din <= 32'h73368775;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07e; din <= 32'h31d35c9c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00b; din <= 32'h0e5ee083;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h356; din <= 32'heb4573c4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c3; din <= 32'h7cf1b7e5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h246; din <= 32'hf32bc6e5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h036; din <= 32'h691db8fb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h142; din <= 32'h76a01a5a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3de; din <= 32'h02838ade;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h272; din <= 32'h77492f10;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h387; din <= 32'h1e27f8ec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h371; din <= 32'h7e165b3e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b4; din <= 32'h10bb7df7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01b; din <= 32'h87734db3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h240; din <= 32'hc05e9574;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b2; din <= 32'he580b7a8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h278; din <= 32'h932088f1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cc; din <= 32'h66d288cc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b5; din <= 32'haff36a16;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d8; din <= 32'h719ab759;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c8; din <= 32'h5f87c334;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f6; din <= 32'h4ab3c93f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08b; din <= 32'hf64235a2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a3; din <= 32'hd8aa74e1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f2; din <= 32'hd0fe90e9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h073; din <= 32'hf2316f61;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ee; din <= 32'h8c2993c3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h106; din <= 32'h6035b954;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h209; din <= 32'h68fc54ba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24e; din <= 32'h634b7f66;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2af; din <= 32'hb90ee4dc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h294; din <= 32'h765dfb2a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c8; din <= 32'h02db7fb9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h029; din <= 32'h038904e9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b4; din <= 32'hfd8d7ae0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h200; din <= 32'hfe0415cf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c8; din <= 32'h3df89ae5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29e; din <= 32'hd559b5e7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00b; din <= 32'h83873f64;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f0; din <= 32'h3b37c995;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c6; din <= 32'hf11fb744;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ea; din <= 32'h92f17e77;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h293; din <= 32'h5a610cbb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b2; din <= 32'h7df04d98;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h115; din <= 32'h8ae0e702;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bd; din <= 32'h8b632acc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h391; din <= 32'h96a0897c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fd; din <= 32'hc4a541be;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e1; din <= 32'hf2d4762e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h388; din <= 32'h57b542b0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c2; din <= 32'h7b43a63c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f9; din <= 32'h1c54e9bc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f1; din <= 32'h6768cd67;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h390; din <= 32'hb2f1f22a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22c; din <= 32'h272bf83f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d2; din <= 32'hb31dfbd7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27e; din <= 32'h4210f94e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h369; din <= 32'he042db31;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bd; din <= 32'h0cdb8f59;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h017; din <= 32'h0a4e6fa3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e6; din <= 32'h3c49ec27;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ca; din <= 32'h5bbb98a4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e9; din <= 32'h5914c461;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h212; din <= 32'hba092e75;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d9; din <= 32'h11f48f94;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23f; din <= 32'h321757ed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36f; din <= 32'h46dbf78a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d0; din <= 32'h4c14a6dc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h387; din <= 32'hbe4490f7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h219; din <= 32'hee011a83;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13c; din <= 32'h0e095ce1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b8; din <= 32'h6aa0cb48;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h124; din <= 32'habeaa23e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ab; din <= 32'h9e9f1366;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h325; din <= 32'h250f722c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e3; din <= 32'h74033bcc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h219; din <= 32'hfd8c88fd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h196; din <= 32'hce2a716a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h103; din <= 32'h48041c6b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h275; din <= 32'haeb2fe3d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h379; din <= 32'h6b173b14;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h256; din <= 32'hbddfb16a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h074; din <= 32'h6353a3d3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d7; din <= 32'h9769f3a5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c6; din <= 32'hb211373f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h372; din <= 32'h89489b05;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h098; din <= 32'ha78730e4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h161; din <= 32'h05778d0d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12f; din <= 32'h0b0fbf32;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c5; din <= 32'h4476a4a5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h079; din <= 32'h46205d21;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h336; din <= 32'hc561e130;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bb; din <= 32'hd69aaaa2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h214; din <= 32'hd076235c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d1; din <= 32'he7df1eb7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0dd; din <= 32'hffab151c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03d; din <= 32'hd3c8636b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h140; din <= 32'hfe89d72d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h123; din <= 32'h263dbb87;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h360; din <= 32'h05798751;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h363; din <= 32'h20013ade;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b5; din <= 32'ha5ddb421;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25e; din <= 32'hc9d25145;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38f; din <= 32'h51585883;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b6; din <= 32'h02a1d24f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h163; din <= 32'hbfe53a34;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1de; din <= 32'h2cf3c362;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25d; din <= 32'h20fa4af9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10c; din <= 32'h6e1cd204;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21e; din <= 32'h973f7e9c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h100; din <= 32'h5d7c72ec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bb; din <= 32'hefd944b8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22b; din <= 32'hadb69e50;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e4; din <= 32'h27e20ce5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h156; din <= 32'h341e3c09;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h005; din <= 32'h649177bf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h054; din <= 32'h635e202f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e9; din <= 32'h762b9cf3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a8; din <= 32'h1a0badc1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h200; din <= 32'h866de36b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13f; din <= 32'h7489b231;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e4; din <= 32'hb18c4f33;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f0; din <= 32'h213c975e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f6; din <= 32'h0b90c51c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h136; din <= 32'ha9dac2db;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h279; din <= 32'h8627258f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11c; din <= 32'h3967966b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0aa; din <= 32'h3792688d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36a; din <= 32'h9d9055a7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23a; din <= 32'hc391a897;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24c; din <= 32'h217124ca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c5; din <= 32'h579c7bf3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a6; din <= 32'hc7235627;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31a; din <= 32'hca899b44;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h069; din <= 32'h63bad3f4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e9; din <= 32'he4c4b177;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cf; din <= 32'hf2bfa9e9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h310; din <= 32'h539c645c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h217; din <= 32'h6eb91377;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h263; din <= 32'h5d1a86d9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h240; din <= 32'ha1794ffa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h355; din <= 32'ha6fe85ff;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01a; din <= 32'hd2c59f62;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h165; din <= 32'he367fb36;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h237; din <= 32'h4c14b28b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h042; din <= 32'hb003588b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h086; din <= 32'hb4aa8909;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01c; din <= 32'hc086e727;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2fc; din <= 32'h0a9cda07;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f1; din <= 32'hdfc805d7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ac; din <= 32'h22a44f87;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08e; din <= 32'h094b0c51;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d8; din <= 32'hce4c209b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16b; din <= 32'h374e68b6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14e; din <= 32'h66c9bc42;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cf; din <= 32'hc69aeb72;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23d; din <= 32'h1c849fe8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28d; din <= 32'hdbc0de7b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30f; din <= 32'hf5b207f8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h291; din <= 32'h2b3b3f85;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25b; din <= 32'h1c38fec0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h033; din <= 32'h582c6412;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h288; din <= 32'h82f2dd69;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ff; din <= 32'h571646cd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h092; din <= 32'h9a274af8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h342; din <= 32'h11201a59;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b2; din <= 32'h43d950d0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h299; din <= 32'hb55a6a70;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h358; din <= 32'h1f645201;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ad; din <= 32'h24a6b704;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c2; din <= 32'h602c91a5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b9; din <= 32'h7fac7326;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h160; din <= 32'h04d90323;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h012; din <= 32'h9fde945e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h250; din <= 32'h73c2be9b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ae; din <= 32'h2bf18324;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cf; din <= 32'hb5e83f75;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3df; din <= 32'hcd05e626;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h001; din <= 32'h4f9e1640;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09d; din <= 32'hdf11439f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35e; din <= 32'haf1a681e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h242; din <= 32'hd514de12;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f7; din <= 32'hf7cae43c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37e; din <= 32'h62ee0749;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h083; din <= 32'h2cd852b4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h085; din <= 32'hd6b9e9ce;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fe; din <= 32'hf1b0c004;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c6; din <= 32'hddf0375c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h094; din <= 32'h913790ae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h072; din <= 32'h3e229121;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e8; din <= 32'h7ac990ac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27e; din <= 32'hc8f97b6d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09b; din <= 32'hb058baa2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h039; din <= 32'h74016893;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17c; din <= 32'h90384240;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16c; din <= 32'h276cd9a7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h319; din <= 32'hf82fd00f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27e; din <= 32'h8b60bb31;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c9; din <= 32'h90c47c05;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h264; din <= 32'h3429ffec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h250; din <= 32'hbed7aa54;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bb; din <= 32'hb97d394a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d1; din <= 32'h5b9fe1a7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c3; din <= 32'h0fb0dcca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05e; din <= 32'h39e556a5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h389; din <= 32'h0bd497c2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d5; din <= 32'hdfc097b8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h224; din <= 32'hf1dee211;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h100; din <= 32'h6b5a4f5a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ca; din <= 32'hee94efc4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d1; din <= 32'h2e93b789;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a6; din <= 32'h4933c674;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13f; din <= 32'h3b4494a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08e; din <= 32'hc090e710;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01a; din <= 32'hb6f0b45c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h205; din <= 32'h51d8468e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2fb; din <= 32'h7727d782;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1aa; din <= 32'h43da2153;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h103; din <= 32'h5604199a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h041; din <= 32'ha633f003;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h354; din <= 32'h5194745a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00e; din <= 32'h3a91f79c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h364; din <= 32'h624bcd69;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f7; din <= 32'h9fd8d5c4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11d; din <= 32'hc1102c96;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h308; din <= 32'h62c2ae1c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e4; din <= 32'h6e7664fc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h142; din <= 32'h97a5e98c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h153; din <= 32'h1137c515;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e1; din <= 32'h0c93da72;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28c; din <= 32'h3c9fa038;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h141; din <= 32'h3219989a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16b; din <= 32'hc3973dd5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h182; din <= 32'h8e0fc3ed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bb; din <= 32'h583633bd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h059; din <= 32'ha1c80bcf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ee; din <= 32'h0a8feca4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h303; din <= 32'h1c4f0879;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h045; din <= 32'ha32d039c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c9; din <= 32'h2c45e947;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c2; din <= 32'ha02e01db;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h338; din <= 32'h8a6dd07d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h035; din <= 32'h49c2070c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f5; din <= 32'h20e2fe6a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c1; din <= 32'hd4b68f4d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h272; din <= 32'h9bbf016b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26e; din <= 32'h3c1d7112;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h040; din <= 32'hdcb98e6f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h017; din <= 32'h1aaf1354;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h279; din <= 32'h2f6b55f8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38b; din <= 32'he11298d5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h391; din <= 32'h8be9b69c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a1; din <= 32'hae2bf834;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h156; din <= 32'haec11a0a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h290; din <= 32'h255ff60a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b9; din <= 32'hac4d6ec3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h387; din <= 32'h208c5392;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e4; din <= 32'h93e8aa7d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h008; din <= 32'hb83db0f8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h170; din <= 32'hdd1de3de;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12a; din <= 32'h5fdd2e4f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e7; din <= 32'hcc01bd67;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h297; din <= 32'hf1be9723;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h026; din <= 32'h42950ee0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14b; din <= 32'h79e4bfef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ca; din <= 32'h8fef85cc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h255; din <= 32'h9390923a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h324; din <= 32'h100d757e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13a; din <= 32'h48ffdf44;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h067; din <= 32'h4a2cf483;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3be; din <= 32'hfd545aef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h199; din <= 32'h2958915b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f0; din <= 32'hca17ea50;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a4; din <= 32'hf877636e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h059; din <= 32'ha8373186;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a9; din <= 32'ha2b12d1d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h346; din <= 32'h01b44e5f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36f; din <= 32'he3dbb075;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h226; din <= 32'ha8b03298;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b3; din <= 32'h1fb87d02;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ac; din <= 32'h1e6be0a4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a3; din <= 32'h59b5a27a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ff; din <= 32'h984cc725;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fa; din <= 32'hc1e6e6ad;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h024; din <= 32'hba428366;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05e; din <= 32'he63919c2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04e; din <= 32'hadcdcccd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h337; din <= 32'hb10b1447;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c1; din <= 32'hd0efa821;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cd; din <= 32'h29f9e39a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f5; din <= 32'hf1f8b53a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h238; din <= 32'hce90f0af;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h352; din <= 32'h3f7a7331;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h367; din <= 32'h678436e9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h193; din <= 32'h82939f22;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c1; din <= 32'h7c534b71;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36d; din <= 32'ha4cfe772;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h142; din <= 32'hcef4dfaf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h354; din <= 32'h652e7652;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h255; din <= 32'hb1c2d88b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h216; din <= 32'h382591b2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h230; din <= 32'h9db7512a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h218; din <= 32'ha30dfb29;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h047; din <= 32'h3ea54e71;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h369; din <= 32'h3f1113a8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f2; din <= 32'h27878dd1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h145; din <= 32'hc85a5442;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2dc; din <= 32'h9ed8c53e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h105; din <= 32'h7135e598;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3dc; din <= 32'hd91ecb9b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d2; din <= 32'hc7366a0f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e8; din <= 32'hff98b992;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d7; din <= 32'h776c085e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h140; din <= 32'h74e3e8bb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b1; din <= 32'h8eea41d4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b5; din <= 32'hf298aead;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h326; din <= 32'h15ad450d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06f; din <= 32'h421266da;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31c; din <= 32'h77546746;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c7; din <= 32'h76276eba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h329; din <= 32'h35be6b80;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h222; din <= 32'h266b91eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h292; din <= 32'h6c670b67;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1de; din <= 32'hc9a455de;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h082; din <= 32'hc64fd8ee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e4; din <= 32'h41a1f97c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bf; din <= 32'hfab81d7a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ce; din <= 32'h2476c499;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h069; din <= 32'h9d73a5ce;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h067; din <= 32'h1ccc3f95;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f1; din <= 32'hc0a5a18e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28a; din <= 32'h5da8ac84;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h096; din <= 32'h6d4a27ae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f9; din <= 32'h87708e2b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h124; din <= 32'ha542ecaf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d3; din <= 32'h38ee3825;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h001; din <= 32'hb73d83af;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07a; din <= 32'hda1ca887;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35b; din <= 32'h85b4e589;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b5; din <= 32'hc7c52e93;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f4; din <= 32'hbb3bf2c5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39f; din <= 32'h94d0809f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h305; din <= 32'habc08e19;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f4; din <= 32'h2c6cd4e9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c8; din <= 32'hb9c39678;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28d; din <= 32'hc8f7783d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2af; din <= 32'hcccc9238;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a8; din <= 32'h8083fcd1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d6; din <= 32'hf7870340;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h185; din <= 32'h50f69c80;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cd; din <= 32'h99110d27;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c0; din <= 32'h7e5315c5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b8; din <= 32'h40f669b5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26c; din <= 32'h89ce20b0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bb; din <= 32'h4f9a0ecb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a2; din <= 32'hf384a323;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h264; din <= 32'he46908c0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b8; din <= 32'he85dfc24;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b2; din <= 32'hcc38a70f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b6; din <= 32'h4e372875;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bf; din <= 32'hd5858d0b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06c; din <= 32'h6d96f747;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16f; din <= 32'hb4b68528;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h027; din <= 32'haacc1b63;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h061; din <= 32'h7244ba82;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f9; din <= 32'h5f9bdbde;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01c; din <= 32'h8ad5af1d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h066; din <= 32'h85d5a864;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13b; din <= 32'ha5604e8a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h139; din <= 32'hef16ebe2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d0; din <= 32'h11bbefc0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h372; din <= 32'h2b4f6041;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h225; din <= 32'hf09993b0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h209; din <= 32'h030d31ff;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f1; din <= 32'hbdbab95a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32d; din <= 32'h14d77d54;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37c; din <= 32'h9c17e2df;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28b; din <= 32'hd5c6a4c6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a2; din <= 32'hfe8493fe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a4; din <= 32'h7ad0347a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b1; din <= 32'h1e5f5a83;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00e; din <= 32'h38dc8852;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h155; din <= 32'h1fdf0025;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e4; din <= 32'he99b4ff9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15b; din <= 32'h37320c1b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h226; din <= 32'hac81e5bd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b8; din <= 32'h19f6bdb7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33a; din <= 32'h93a2fdbc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h025; din <= 32'h781ff7dd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h209; din <= 32'hffba1977;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h055; din <= 32'h3bd631e4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c0; din <= 32'h9c70873c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01b; din <= 32'hb408f586;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h124; din <= 32'h30901800;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h140; din <= 32'h3fcf87e9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fe; din <= 32'hd316b159;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ac; din <= 32'hfdbcd4e7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02f; din <= 32'h5d4a4d9a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h060; din <= 32'hede44f78;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h276; din <= 32'hc09906df;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h018; din <= 32'ha23b0aa0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07f; din <= 32'h70b6e13f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h276; din <= 32'h5ce8a767;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h171; din <= 32'he672785e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20d; din <= 32'h45062438;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28b; din <= 32'h12c67a9b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h227; din <= 32'hd7a9efac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02c; din <= 32'hc311bd3e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h306; din <= 32'hd12a82d2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h014; din <= 32'h4680689e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h165; din <= 32'hec11a71c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h269; din <= 32'h42ab1feb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f1; din <= 32'h8ab8b7c4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f8; din <= 32'hd1173b5b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e5; din <= 32'h146c810f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h384; din <= 32'hb2c98fbd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cd; din <= 32'he4093e28;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ef; din <= 32'h4c2b0c16;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c9; din <= 32'h3bd4c869;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26c; din <= 32'h68421a6b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2af; din <= 32'h96063aaf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h277; din <= 32'h17d6ae20;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h365; din <= 32'h33930a86;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h208; din <= 32'h6239c6b7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h085; din <= 32'h97c6b69d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h361; din <= 32'h07cac535;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h106; din <= 32'hfbeb181b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h280; din <= 32'h223be605;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h048; din <= 32'h318b64bd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23e; din <= 32'hf8390197;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h289; din <= 32'h8a997c47;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h158; din <= 32'hbeb03358;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a0; din <= 32'hfb567476;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17f; din <= 32'hd8605ce9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h177; din <= 32'hb903c482;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26f; din <= 32'hb23e0b4a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h230; din <= 32'h88facecb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0db; din <= 32'ha0d24b9c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e1; din <= 32'h59b69d41;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a7; din <= 32'h8e6ad4fb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h021; din <= 32'h41580372;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06b; din <= 32'h99cc0972;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h019; din <= 32'hbbc6a4ad;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b2; din <= 32'ha61816a2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h231; din <= 32'h791875cb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h217; din <= 32'h786ea4d8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c5; din <= 32'h8eaa1f52;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0de; din <= 32'hf07fa777;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06b; din <= 32'h3bab85a3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h099; din <= 32'h7654e044;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h313; din <= 32'h1f165b7e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3eb; din <= 32'h30201dba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e5; din <= 32'h50a8005b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10d; din <= 32'h01658edb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h283; din <= 32'h3f0de025;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22e; din <= 32'hdcd7fced;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a0; din <= 32'h98046ea2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18c; din <= 32'h6cd11e79;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28b; din <= 32'h1a1cf91a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h350; din <= 32'hcfbbbf13;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fb; din <= 32'h2c634ab4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h069; din <= 32'h6aedfda8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27e; din <= 32'h2f5fc76e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h030; din <= 32'h655cf314;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h372; din <= 32'h6858e872;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30e; din <= 32'h1bf833d4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2df; din <= 32'h8af60295;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d4; din <= 32'h7c3937b8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h368; din <= 32'he719692b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0aa; din <= 32'h53d4142b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f5; din <= 32'hda2d1114;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h352; din <= 32'hdf354cb8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38a; din <= 32'h34715dd8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ae; din <= 32'h111fd24c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24a; din <= 32'hcc902ed1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c0; din <= 32'h9c5b4663;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h032; din <= 32'h5e029ce9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31f; din <= 32'h1df84125;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fa; din <= 32'hbfcaa737;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fb; din <= 32'hfcabca10;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h193; din <= 32'h20f4dfb3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1af; din <= 32'h4a96ac48;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h340; din <= 32'h27899ac3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h398; din <= 32'hd37e0157;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30d; din <= 32'h86d7e330;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h238; din <= 32'h4ea84658;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h285; din <= 32'h3c27412f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h085; din <= 32'h5a655d1a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b7; din <= 32'h93c35ade;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h215; din <= 32'h0cf49748;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cf; din <= 32'hfd3dcb79;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d8; din <= 32'h8952f7fc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h005; din <= 32'h63a78260;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h255; din <= 32'h01ec9d16;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e5; din <= 32'h7e4627b5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13b; din <= 32'ha12cf9ef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08e; din <= 32'h3ab7b8cb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h397; din <= 32'hec1dc377;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a4; din <= 32'h089cac0a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1da; din <= 32'hb2f0051e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c1; din <= 32'h58e19ab6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e2; din <= 32'he8427a1a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h309; din <= 32'h4c7b5278;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h230; din <= 32'h9b05d019;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ae; din <= 32'h3e6c7061;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35e; din <= 32'h9b211106;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e2; din <= 32'hc08f3c31;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30c; din <= 32'h29ca46ef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h247; din <= 32'hfe56fe93;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h022; din <= 32'h33f12c1e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h186; din <= 32'hcd429442;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26d; din <= 32'hb16c50a1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h211; din <= 32'hc278f106;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d0; din <= 32'h0c25b061;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h137; din <= 32'h52b048a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h182; din <= 32'h91f0b0fa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31f; din <= 32'h522844f0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h356; din <= 32'hc093da78;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h215; din <= 32'h8e12bc89;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26b; din <= 32'h394216b6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2db; din <= 32'h8d0d65bf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13c; din <= 32'hc0779f93;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31e; din <= 32'h2e62e345;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00b; din <= 32'h2cf3f0ce;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c8; din <= 32'h32c0a59b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30f; din <= 32'hc760f1ed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ee; din <= 32'he8965e4e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c9; din <= 32'h50b3ceeb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d6; din <= 32'h6f90ee0e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ef; din <= 32'h0fe64c19;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a3; din <= 32'hb73b7c69;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02f; din <= 32'he6f0db15;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25b; din <= 32'h38cefa6d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e0; din <= 32'h04c87462;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h222; din <= 32'h99a2257f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02d; din <= 32'h95024dc7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30f; din <= 32'h670103f2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h322; din <= 32'hb4a6ecec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b1; din <= 32'hb1f7ca56;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c9; din <= 32'h2a3eb454;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h380; din <= 32'ha6fd274a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06b; din <= 32'h23525e59;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c0; din <= 32'heac1672b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0af; din <= 32'h3c86f00f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19f; din <= 32'h96fa223c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38c; din <= 32'hd36adb98;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36d; din <= 32'h6f16c0ed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c7; din <= 32'h553ba355;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b4; din <= 32'ha3484637;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h197; din <= 32'hffe6633f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b9; din <= 32'h83c8e651;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h118; din <= 32'h8a1ffa82;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h366; din <= 32'h5f04c276;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h322; din <= 32'hf0d6b60c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ab; din <= 32'h23a6e631;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h019; din <= 32'h38847c62;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d3; din <= 32'h4f427acc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f4; din <= 32'h8c25a0b9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h169; din <= 32'h4e2126b7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fc; din <= 32'haecbfe5d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h297; din <= 32'h56571080;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26c; din <= 32'h0742751b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h371; din <= 32'h9b62b1a7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h361; din <= 32'h566c921f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30e; din <= 32'h4aae9277;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33c; din <= 32'hb7720986;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h151; din <= 32'h2afcf4eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ed; din <= 32'h916dc991;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2aa; din <= 32'h5ab65328;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22d; din <= 32'hd2d35300;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0af; din <= 32'hc3949a7c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a8; din <= 32'h711fe76a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2fd; din <= 32'hd4f47fce;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h325; din <= 32'h6a22fbb3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ec; din <= 32'hea6b7044;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05e; din <= 32'h52bf9836;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h243; din <= 32'hdc1def09;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h262; din <= 32'hc759ffe8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h214; din <= 32'h8e6f2358;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00e; din <= 32'h3a8c44cb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h210; din <= 32'h6d018e52;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13b; din <= 32'h45567cd3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h157; din <= 32'h26a73809;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30e; din <= 32'hd333ae04;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h005; din <= 32'h33b95c0c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36d; din <= 32'h7289fb14;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e2; din <= 32'h20be765b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c9; din <= 32'h3533fa4f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f2; din <= 32'hdbd621ae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h023; din <= 32'hc0c3c887;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h288; din <= 32'hf90e0f67;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e3; din <= 32'h5bc98355;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39b; din <= 32'hc94233ae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h346; din <= 32'h52ab8da2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17a; din <= 32'h6394f4fe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09f; din <= 32'h6511ac29;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h115; din <= 32'h9e1c3dfc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08b; din <= 32'h09d28edd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13e; din <= 32'h0c50b567;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e0; din <= 32'ha96b2900;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f1; din <= 32'h5ee75f6c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11b; din <= 32'h8ecb13e9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h366; din <= 32'h5485be4d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28a; din <= 32'hf66af26d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h004; din <= 32'he8fe0590;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29e; din <= 32'h3772d857;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h096; din <= 32'h555e1885;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h058; din <= 32'hf4a9743f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20d; din <= 32'h586715b3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28e; din <= 32'hff764d55;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h175; din <= 32'h5e8b902e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ec; din <= 32'h9f0431b6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h350; din <= 32'hb87a96cb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f6; din <= 32'h0f77ce56;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27e; din <= 32'hebced6d3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h273; din <= 32'h056047f0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bd; din <= 32'h23c7144f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h389; din <= 32'h347ccd32;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3dc; din <= 32'h71a61966;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h080; din <= 32'hd3b16046;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h224; din <= 32'h4ef924e2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f3; din <= 32'he968f460;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ed; din <= 32'h259ee023;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ba; din <= 32'h7b085ee2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h049; din <= 32'hf3bb64b9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h020; din <= 32'heb0359c8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14c; din <= 32'habb42497;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h328; din <= 32'h4bde32d9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31b; din <= 32'h3b8767cc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h373; din <= 32'h117a2f07;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16f; din <= 32'h0d3034db;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01a; din <= 32'h674d0096;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c1; din <= 32'h315967eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h375; din <= 32'ha4918728;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3af; din <= 32'he7def603;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h336; din <= 32'h941e18b3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h265; din <= 32'he8654676;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3af; din <= 32'hdbaa7158;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fa; din <= 32'haddcba26;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b7; din <= 32'h752429aa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ee; din <= 32'hf6d59e9e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a6; din <= 32'h50343af6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b4; din <= 32'h4d8ea6aa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34b; din <= 32'h47eb7295;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h277; din <= 32'h546622c2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d6; din <= 32'he858d1ba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12d; din <= 32'hec64d71d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01c; din <= 32'hd8b48ddb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07a; din <= 32'h28cfe0c2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h248; din <= 32'h11071235;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h382; din <= 32'h48beafc1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ac; din <= 32'haf2c353e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13b; din <= 32'h36b9abe9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0dd; din <= 32'h637337a9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06c; din <= 32'hdfd2e55a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04b; din <= 32'h8e9fa761;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2de; din <= 32'hffc04d65;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18c; din <= 32'h65440d11;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02b; din <= 32'h7de66fe3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h159; din <= 32'hae129667;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28e; din <= 32'h0c87d387;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h190; din <= 32'h2751f204;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e4; din <= 32'h5faf2b3b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h149; din <= 32'h43344b20;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h163; din <= 32'h61b7f2aa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b5; din <= 32'hcc6e5309;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ee; din <= 32'h4d565e70;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h080; din <= 32'hbbdb4991;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h110; din <= 32'h6c126c1d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h102; din <= 32'h08ab6132;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h112; din <= 32'h313c6763;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24f; din <= 32'h750750aa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h102; din <= 32'h03140bb6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10e; din <= 32'h5e2e5369;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f1; din <= 32'h07e0a768;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1eb; din <= 32'h38e7ad18;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h120; din <= 32'h7b79823f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h399; din <= 32'h5f0f5634;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a7; din <= 32'h6a03766c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33e; din <= 32'h427079fa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0eb; din <= 32'hddebc893;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2de; din <= 32'h930170df;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fb; din <= 32'h01dbcb50;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h104; din <= 32'h39262e56;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e9; din <= 32'h63ef487c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fa; din <= 32'h180c3c40;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c4; din <= 32'h56dfe52a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h237; din <= 32'h48b59743;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h026; din <= 32'h277a1f76;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07a; din <= 32'he1b0546e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1de; din <= 32'h027bced3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bf; din <= 32'hab0efaf8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h393; din <= 32'h88fdc3c6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h154; din <= 32'hffb03f23;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h219; din <= 32'h9c329bc6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h214; din <= 32'h955ae6b5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35f; din <= 32'h098e2fac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f1; din <= 32'h8cd3f5e3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h375; din <= 32'h7ed10ffa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38d; din <= 32'h438c4dd5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h153; din <= 32'he867adfc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ad; din <= 32'hf53d4cb3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h134; din <= 32'h6b8a733c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ec; din <= 32'h93d4432b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13c; din <= 32'h2f78866e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10e; din <= 32'hc9407c23;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h016; din <= 32'h56e0cd37;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b6; din <= 32'h1db28185;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h258; din <= 32'h9ef31bc4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h386; din <= 32'h0be2c4f5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a6; din <= 32'h74072360;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e1; din <= 32'h7f03230a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f6; din <= 32'ha6aae02a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h127; din <= 32'hd085ca93;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23f; din <= 32'ha62e7f28;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e9; din <= 32'h8cf92891;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h044; din <= 32'h94e2fd51;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h017; din <= 32'h93bf0223;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h111; din <= 32'h2b422d86;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h352; din <= 32'hcefa49af;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0eb; din <= 32'h823f441d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10e; din <= 32'h64fd069d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h263; din <= 32'h4f2513f5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f7; din <= 32'h0dcb9a2b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c8; din <= 32'h3e0a62a5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h236; din <= 32'h640811b0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32d; din <= 32'h03f56a07;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h318; din <= 32'ha52b68c8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16e; din <= 32'hd820cf03;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h083; din <= 32'hae73111d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h016; din <= 32'hff526304;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bf; din <= 32'hd48d99a9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05e; din <= 32'h971d8d4c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d9; din <= 32'h6b5f5d0b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f3; din <= 32'h8d019077;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a1; din <= 32'hed1600b4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22e; din <= 32'h3919a899;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15d; din <= 32'h821a8b3f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h376; din <= 32'haeea5f26;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h234; din <= 32'h5bc099b9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f1; din <= 32'hc4b4598a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h216; din <= 32'h02aa3239;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h298; din <= 32'he74a1649;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36a; din <= 32'ha4d45581;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31c; din <= 32'h75d7bbdd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ea; din <= 32'h9a80b0c2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e1; din <= 32'hdaaa4b4b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h010; din <= 32'h44d8bb9e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c5; din <= 32'h32741dde;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d5; din <= 32'hc9edba07;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h107; din <= 32'h172bde61;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f1; din <= 32'hc061bdb4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h303; din <= 32'h44068bad;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a6; din <= 32'ha7a82b0f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h214; din <= 32'haa1cba0f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1aa; din <= 32'h24f63539;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h145; din <= 32'hdee7e00e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28c; din <= 32'hfb45b231;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h195; din <= 32'h79d173f2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cb; din <= 32'h47c0ea23;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h001; din <= 32'h3d2c4c97;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e3; din <= 32'h9b386c58;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3da; din <= 32'h1956868b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e9; din <= 32'h2d5933db;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h063; din <= 32'he6b66abb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h380; din <= 32'h821091b4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13c; din <= 32'h21e38768;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h028; din <= 32'h6493793b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f8; din <= 32'h6fdadac0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f0; din <= 32'hdec3a359;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24e; din <= 32'h37f782c9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28d; din <= 32'hb9a81f06;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22e; din <= 32'hf1eaa2c3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h295; din <= 32'h3d4cfc83;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b7; din <= 32'h32f09757;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b9; din <= 32'h8278328f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e0; din <= 32'h91a49fc3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29f; din <= 32'h10bd25f9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h233; din <= 32'h3f91bef6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12c; din <= 32'hc9c1037b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h342; din <= 32'hea834bf5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14d; din <= 32'hd949d56f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12a; din <= 32'hf1d9060c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e6; din <= 32'h111548c6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2db; din <= 32'h7abc7dde;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b8; din <= 32'h3297faf5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00c; din <= 32'h9deb072d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30b; din <= 32'h426d827e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h057; din <= 32'h21cdfd94;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f7; din <= 32'hc6b3dd9a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14e; din <= 32'hcaf2e8f0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h102; din <= 32'h3bd8cdc6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f6; din <= 32'hfdc28b47;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b8; din <= 32'hbe79ff06;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f2; din <= 32'hefb5bdbf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b7; din <= 32'hfc42d239;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33e; din <= 32'hc3e45045;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h317; din <= 32'h6c6183e3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h339; din <= 32'h1e2a4bde;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30a; din <= 32'hc81fadde;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ba; din <= 32'h0b591a6c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e8; din <= 32'h6d2dda03;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a3; din <= 32'h95160e0e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fb; din <= 32'hd3a63478;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29a; din <= 32'h9d64fcb6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h267; din <= 32'hc85adb5f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h021; din <= 32'he0efbbfe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30f; din <= 32'hf68aff5e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15e; din <= 32'h8652985c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03a; din <= 32'h3eacfa19;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h046; din <= 32'hecd950f6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e3; din <= 32'he98b06dd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2eb; din <= 32'h5475ad8d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h277; din <= 32'hf83a3eb1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h190; din <= 32'h4ff03f38;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d7; din <= 32'h25610ea6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h293; din <= 32'hfdfbd674;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h057; din <= 32'h458e4fc2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c6; din <= 32'h0405b7b2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h316; din <= 32'h265311a2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f9; din <= 32'h28066f41;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b3; din <= 32'hb73e13ae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c1; din <= 32'hea8fd3ba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e6; din <= 32'h64586dcc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14a; din <= 32'h1958edb1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h319; din <= 32'h07d132ff;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e9; din <= 32'hcf754c8a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e2; din <= 32'haf191743;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h339; din <= 32'hdfc776e5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h209; din <= 32'h3073fc82;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25b; din <= 32'h63fdfe5e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cb; din <= 32'h0a10303e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32d; din <= 32'hdbd3cf22;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h354; din <= 32'h67e2a57f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c8; din <= 32'h6edceb49;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3eb; din <= 32'h1e9fced2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e4; din <= 32'hbbf9257b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16e; din <= 32'h9774435e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h202; din <= 32'hd012395b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20d; din <= 32'h5040d6ce;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c3; din <= 32'haf5d953f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h376; din <= 32'h19d430ef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e3; din <= 32'h2b3d8c28;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09d; din <= 32'hecb0980b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ee; din <= 32'hae530352;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h156; din <= 32'h42a733ea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b7; din <= 32'h3ae79233;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10c; din <= 32'h87f08db0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e4; din <= 32'h235e1a9a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0af; din <= 32'hd647fc68;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f4; din <= 32'hf41b7d9e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2dd; din <= 32'h3c6c8a92;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ec; din <= 32'hce044bb7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0be; din <= 32'h4844eb3f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h394; din <= 32'h810f4952;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02a; din <= 32'h8c5db6d8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17a; din <= 32'he1c648bd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f6; din <= 32'hd65f2710;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26e; din <= 32'h37cbfe36;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32e; din <= 32'h198b3afa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d8; din <= 32'h94df7ee9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b5; din <= 32'h65d0d9fa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38f; din <= 32'h136cc56e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31b; din <= 32'h9435cf8f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h365; din <= 32'hb5ad68fe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20d; din <= 32'h44bd3fc3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e3; din <= 32'hb3267884;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h208; din <= 32'hd81caa19;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c9; din <= 32'h1454b0c1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h009; din <= 32'h5529f07d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h327; din <= 32'h8639801e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18f; din <= 32'h577ddf7e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h141; din <= 32'he5094922;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14d; din <= 32'h6cee2698;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h158; din <= 32'hc9045054;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a9; din <= 32'hdf0d9e69;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29f; din <= 32'hdb6ddfba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b5; din <= 32'h1e5ee4b6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h081; din <= 32'h5f44e633;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b7; din <= 32'haa0b5591;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h305; din <= 32'hf09fa2d9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3db; din <= 32'hec3d6dcd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a1; din <= 32'hc4e7c786;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h205; din <= 32'hf0a14188;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c6; din <= 32'h8db440ae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h129; din <= 32'hca742351;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b4; din <= 32'h910adf57;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h011; din <= 32'hdb90f54c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h244; din <= 32'h5ec037ef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h208; din <= 32'h2ac258a7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23b; din <= 32'h8c8ca90c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h373; din <= 32'h307eb4a5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2df; din <= 32'hecafad79;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h240; din <= 32'ha521422a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ca; din <= 32'h8a5253b5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37e; din <= 32'h2081950e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c8; din <= 32'h857b45cb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2dd; din <= 32'hdf5c2fff;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ab; din <= 32'hc4b32717;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ee; din <= 32'he2161386;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h218; din <= 32'h1f8df8a3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h016; din <= 32'h775583e7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h353; din <= 32'he6b3b847;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fa; din <= 32'h735f9aa3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28e; din <= 32'h1bc4d8f0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h213; din <= 32'hf9a43af2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h024; din <= 32'h482b8d91;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12a; din <= 32'hb4edfddb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h373; din <= 32'hc2af1cfa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37c; din <= 32'h3f988d86;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12f; din <= 32'h50fa1283;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h236; din <= 32'h8fdc979a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h252; din <= 32'hc947b369;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h198; din <= 32'h82517d2a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h126; din <= 32'h4e7d5f2e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c7; din <= 32'hb5b42e80;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26e; din <= 32'h4c678415;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ed; din <= 32'h0dc5878b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h222; din <= 32'h579a78b4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25a; din <= 32'hc8c1b11e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e5; din <= 32'h62a3e14a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fe; din <= 32'h1a6951aa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e1; din <= 32'h6dcd9651;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h046; din <= 32'he9ec5209;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38d; din <= 32'h808e150e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bc; din <= 32'hff985cc7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ac; din <= 32'he0da3047;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h087; din <= 32'hbd166106;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h118; din <= 32'h698a40ed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bf; din <= 32'h4ce7c247;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03f; din <= 32'hce070c45;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cf; din <= 32'h70bb999c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h073; din <= 32'h3838f80d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02b; din <= 32'h5b6d11c5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f5; din <= 32'h36d6b15b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h206; din <= 32'hbc0a395c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3af; din <= 32'h6d75bfd8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h335; din <= 32'hb2885555;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00c; din <= 32'hda4c1328;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02a; din <= 32'h0bf56c3f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e8; din <= 32'hc0166daa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e2; din <= 32'hec1b1c32;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a8; din <= 32'h24837301;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h007; din <= 32'hf1e56e5f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e1; din <= 32'h46fef419;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h360; din <= 32'h0529d683;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cf; din <= 32'h51e684a9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c8; din <= 32'h594b6afa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h296; din <= 32'h3e4098c7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c2; din <= 32'h7a2dfa0a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h382; din <= 32'hf05b5124;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d4; din <= 32'hcec3d5c4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d7; din <= 32'hb4004fea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cf; din <= 32'hb377f1b0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cc; din <= 32'hdb2c7b79;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24e; din <= 32'h8877ce1f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d3; din <= 32'hf48f746c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e1; din <= 32'h9d130da9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b3; din <= 32'h41221957;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13e; din <= 32'h7e5bcf2a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h133; din <= 32'hbddef7d9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32d; din <= 32'hcf40d1a4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34c; din <= 32'h2ca68e04;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f0; din <= 32'h448b51ff;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h184; din <= 32'hda4ea896;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22b; din <= 32'hb8693e84;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h339; din <= 32'hda39e1a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c3; din <= 32'hd7cd8926;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3dd; din <= 32'h9764f0e5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37b; din <= 32'h661f756c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20e; din <= 32'heef9ba8b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cf; din <= 32'hfccd4039;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h245; din <= 32'h114a230a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h001; din <= 32'h69aaba61;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14d; din <= 32'hc65ed78d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14f; din <= 32'h15fb2536;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h269; din <= 32'hb0c102e0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17f; din <= 32'h4fa0f449;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17d; din <= 32'h0b63682d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ca; din <= 32'h3e34e7ef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h185; din <= 32'h28471cb5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f3; din <= 32'h01981099;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ac; din <= 32'hc60bcab8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h304; din <= 32'h001a26a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b1; din <= 32'h9d67b6ab;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f7; din <= 32'ha8b20f2b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h259; din <= 32'hcceb103b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fc; din <= 32'h24a3707c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h317; din <= 32'he975aca0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bc; din <= 32'hdbad6fa4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b7; din <= 32'hd6cccb85;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ad; din <= 32'h8c14b83c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ce; din <= 32'hf43fb711;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29b; din <= 32'hb21288be;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a4; din <= 32'h64ecb70a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cf; din <= 32'h296586a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d5; din <= 32'h4c88cbf6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c0; din <= 32'h5fce7b9f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2db; din <= 32'h153c9459;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21d; din <= 32'h28bb4d0d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h354; din <= 32'he54f9dd2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h363; din <= 32'h44635b83;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34b; din <= 32'hcf0a3b63;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27a; din <= 32'h59befe69;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d2; din <= 32'h62da238b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h017; din <= 32'h6b7497d5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h212; din <= 32'hee2fec8b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ba; din <= 32'h1b639fcd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d4; din <= 32'ha1b61692;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20f; din <= 32'hd6326818;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fc; din <= 32'h67a114f4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h133; din <= 32'h908af57f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b9; din <= 32'hf961a98e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h246; din <= 32'h3fdeaa5e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d8; din <= 32'he87be84b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31a; din <= 32'h559659a7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h081; din <= 32'hae33e4a7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h258; din <= 32'h6f104b14;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a0; din <= 32'ha9791a91;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h024; din <= 32'h16d531bc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h363; din <= 32'h0c59072c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h327; din <= 32'h571fa712;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h128; din <= 32'h737ad8aa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ef; din <= 32'he52d7df2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h181; din <= 32'hd9f0ecc3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h309; din <= 32'hfcfa78b1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f6; din <= 32'hb3fcf619;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22e; din <= 32'hd1003715;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37d; din <= 32'h5c33df3c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3dd; din <= 32'h260afc97;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h181; din <= 32'hfb11843a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cb; din <= 32'hc25aac85;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29e; din <= 32'h08b8b0dc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h296; din <= 32'h6b8015aa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38a; din <= 32'h3f9f107e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h045; din <= 32'he0d6aea3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24d; din <= 32'ha62aacc7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h102; din <= 32'hd6e875c9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d1; din <= 32'h141012c1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f7; din <= 32'h1c82fb05;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e5; din <= 32'h9c564a99;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h048; din <= 32'h2378ac12;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h144; din <= 32'hfc11fb48;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d4; din <= 32'h2ef96db7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h291; din <= 32'hd3839333;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h368; din <= 32'hee036a10;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h289; din <= 32'hdcf63ec9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26e; din <= 32'hcf21c73a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d3; din <= 32'h51353492;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h276; din <= 32'h0315ad81;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cd; din <= 32'h1966b14a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h005; din <= 32'h7f290ba2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fc; din <= 32'hba5582e0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h159; din <= 32'h18d2cc1e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19f; din <= 32'h95a8791f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h219; din <= 32'h3ed93800;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b1; din <= 32'h8686f921;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h188; din <= 32'h172fed59;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36c; din <= 32'h7948b834;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09d; din <= 32'h43cb02d2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h230; din <= 32'h580485e9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31b; din <= 32'h62855ec5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3db; din <= 32'h021c8d88;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f7; din <= 32'hac6056dc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ab; din <= 32'h4a83fb52;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h094; din <= 32'hb95f9e15;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f4; din <= 32'hdd441c1a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a9; din <= 32'hf6ae6767;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h328; din <= 32'hbaec640f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21c; din <= 32'h973d6bee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25f; din <= 32'h551db229;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e7; din <= 32'h98e597c0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d3; din <= 32'hd4ea8ace;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1af; din <= 32'haba74052;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a0; din <= 32'hae3d3035;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20c; din <= 32'h51eaef12;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h008; din <= 32'h3009524e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ca; din <= 32'h12abd86c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a8; din <= 32'h8116252d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a8; din <= 32'h6c887446;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03a; din <= 32'h482bd12e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04f; din <= 32'hb1b19138;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h071; din <= 32'hda9d2394;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32c; din <= 32'ha2a32e62;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24f; din <= 32'h7efa37ea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h101; din <= 32'hda5068de;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13d; din <= 32'he493636f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h185; din <= 32'h775b9684;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h362; din <= 32'h017d47f7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h278; din <= 32'hce511746;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h243; din <= 32'h6f5cde0d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b3; din <= 32'hf5156442;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h342; din <= 32'h3a84c717;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08d; din <= 32'h20c8bc84;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d7; din <= 32'h98f224fe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e8; din <= 32'ha81cee54;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h355; din <= 32'h883e171d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14e; din <= 32'h2785734c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a3; din <= 32'h847592bf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h167; din <= 32'h8cb5dd3f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f2; din <= 32'hdf7dd52d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h216; din <= 32'haa78e3a8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f1; din <= 32'h5249c55a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h267; din <= 32'hc505face;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h051; din <= 32'he70b1269;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34c; din <= 32'hf5e84b70;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33c; din <= 32'h28111387;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h138; din <= 32'h79fd73bd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ba; din <= 32'hc7514c30;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h086; din <= 32'h46b5f72c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h216; din <= 32'h40ae1379;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07f; din <= 32'h6562360b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ad; din <= 32'hfaca785f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h184; din <= 32'h548f3b00;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e5; din <= 32'hd19a9e9f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fc; din <= 32'hcd8d7e9d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e3; din <= 32'h4797767c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h184; din <= 32'haff31b23;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h196; din <= 32'hcaf3e48e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h110; din <= 32'he5c4e2ba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b2; din <= 32'h269331e0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bd; din <= 32'h9fd75eb8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a5; din <= 32'hbbe4f87c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h371; din <= 32'h97778762;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e8; din <= 32'h7345c520;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d5; din <= 32'h42e2f18c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h148; din <= 32'hc751fb3a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h390; din <= 32'h4826ba93;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b4; din <= 32'h7653d59c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h021; din <= 32'hcf603749;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27b; din <= 32'h0735f28d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bc; din <= 32'h5de9c6c6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h321; din <= 32'h12b37fc1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h260; din <= 32'hfccf67a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a7; din <= 32'hd0628c88;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h180; din <= 32'h8af3af85;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ee; din <= 32'hf7863cd4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h398; din <= 32'h335da5e0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h044; din <= 32'h38a857a5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h291; din <= 32'h922618e0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b2; din <= 32'hf4bd7390;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h210; din <= 32'h00399d39;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h125; din <= 32'h42affa5d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15d; din <= 32'h0ce17ab5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h026; din <= 32'h6bb00fc9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ea; din <= 32'h5810566c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h012; din <= 32'h7f7d9185;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08f; din <= 32'hcda57c0e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1dc; din <= 32'hf01ff4d4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cb; din <= 32'h3f483746;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h256; din <= 32'h1d05098b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ae; din <= 32'hc6dfc26b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e1; din <= 32'h3fc3955f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c9; din <= 32'h0e247a81;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h329; din <= 32'h1dfad722;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30a; din <= 32'h5be02f76;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39a; din <= 32'h6070a878;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fc; din <= 32'h0a79c3e4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h280; din <= 32'hafa68b7b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h210; din <= 32'h523d0d86;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h233; din <= 32'hd31d1696;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h385; din <= 32'h782d6481;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h018; din <= 32'h7b76b779;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h188; din <= 32'hec9decc2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h103; din <= 32'h301c27aa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cc; din <= 32'h5a657e1e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06b; din <= 32'h940a2143;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07d; din <= 32'hc8b67285;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10e; din <= 32'h945cd4ae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e5; din <= 32'he6a7e8a2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bc; din <= 32'h5b20114b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23b; din <= 32'h6549fc38;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c9; din <= 32'ha94bb6fa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h008; din <= 32'h0f162eca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36b; din <= 32'h9db88134;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f0; din <= 32'hecab1495;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36d; din <= 32'ha6b1a3a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h050; din <= 32'hffc7bb0a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h069; din <= 32'hc69d8e6f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h098; din <= 32'h551d48ec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f2; din <= 32'hd5e7d0a7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04d; din <= 32'h371944c1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d3; din <= 32'h13704382;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e3; din <= 32'h08fffc31;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h109; din <= 32'h9703861f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b7; din <= 32'h29b2850f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h226; din <= 32'he42cbf7e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h380; din <= 32'h8286b752;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h183; din <= 32'h34dc6c84;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33c; din <= 32'h30736b1e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h359; din <= 32'hd090ff45;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h386; din <= 32'hae1dd0fb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h097; din <= 32'hf1932045;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ef; din <= 32'h43b94db0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e4; din <= 32'he2027924;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f0; din <= 32'hc371aee6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h035; din <= 32'hb7517964;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h054; din <= 32'h441dda80;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02f; din <= 32'h72d752be;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h288; din <= 32'h0a4b10f2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e4; din <= 32'hd439d18e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a8; din <= 32'h0c491252;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19f; din <= 32'h43646881;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h299; din <= 32'h3e2bf862;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h333; din <= 32'hfc5ad15b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17a; din <= 32'hd26f3682;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f7; din <= 32'h86c1e557;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a9; din <= 32'h55dece71;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36e; din <= 32'hce7bab3e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ba; din <= 32'h83b065b1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a7; din <= 32'h3efd86d5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h131; din <= 32'h567d4373;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25c; din <= 32'h76ebcd79;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f2; din <= 32'h5587b266;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h324; din <= 32'h9205c238;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h204; din <= 32'h2bb349b8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19b; din <= 32'hd66bdccd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39c; din <= 32'h7b95ce57;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h362; din <= 32'h5f715470;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d4; din <= 32'h1a673846;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h085; din <= 32'h9a7800a9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c2; din <= 32'h9f7107e8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h363; din <= 32'h998cb9b3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h173; din <= 32'hb17a2a53;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b5; din <= 32'hc52b1425;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h166; din <= 32'h8967fcbd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h213; din <= 32'hdb4059b9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h239; din <= 32'ha817c4fd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30c; din <= 32'h622a9560;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2eb; din <= 32'h79a82996;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cd; din <= 32'h6e64b23d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d1; din <= 32'hb7edb749;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19c; din <= 32'h7f43f085;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10a; din <= 32'h1590b662;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h141; din <= 32'hb1c223ed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h130; din <= 32'h2f2d8f78;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21a; din <= 32'h24918c4d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h260; din <= 32'h718eb5b8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26e; din <= 32'hbd9f9a15;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33d; din <= 32'h61406893;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h162; din <= 32'h6ebbbc47;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a2; din <= 32'h669cfa7f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h174; din <= 32'h3998bf36;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1da; din <= 32'h0cb33085;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h000; din <= 32'h3fdf57b4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27f; din <= 32'h2341d32b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h092; din <= 32'he57317c8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cb; din <= 32'h149f11a7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h311; din <= 32'h92bd08d9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c8; din <= 32'h681abad9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h133; din <= 32'hbf8d3837;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h399; din <= 32'h4c1f065f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h377; din <= 32'hbeed9fe5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h158; din <= 32'h2cae8027;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f5; din <= 32'hf8fea1b6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h224; din <= 32'h97799188;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18c; din <= 32'h9c3e56d7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2de; din <= 32'hd96cc147;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f7; din <= 32'hace7d434;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h021; din <= 32'h3bd1a42c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h019; din <= 32'h1d6a7c2b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h054; din <= 32'hf96d3f60;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h028; din <= 32'h08989ef7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h067; din <= 32'h12c6f6a3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bb; din <= 32'h78a548f3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h327; din <= 32'h73076c29;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e4; din <= 32'hbfbe2c2f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a4; din <= 32'hfd00f768;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h365; din <= 32'hc9f96c0f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c9; din <= 32'hc9bb777c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h110; din <= 32'hc5d0ab70;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h142; din <= 32'h7d0cb2ed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f3; din <= 32'he1326beb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f8; din <= 32'h808a3410;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33f; din <= 32'h0a36dffc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ab; din <= 32'hd44adaf3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bf; din <= 32'hdb7a2db3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h001; din <= 32'hd881f3ea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h235; din <= 32'h25e23868;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2df; din <= 32'h45b46a1e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c8; din <= 32'h5026b22c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h015; din <= 32'hd4086b1b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cd; din <= 32'h65a7ac21;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h093; din <= 32'h6e3cd1fb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h348; din <= 32'h209a0da3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38b; din <= 32'hd34b4891;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h384; din <= 32'h25737074;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03c; din <= 32'h9468b224;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d7; din <= 32'h469ab421;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h234; din <= 32'h1f38d1cc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a4; din <= 32'he97ba5b2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34e; din <= 32'hcb230eac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12e; din <= 32'h9fd56679;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ea; din <= 32'h9ad406d8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24e; din <= 32'h19a419eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f2; din <= 32'h0a0f3876;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h208; din <= 32'hd6a3b9b4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30e; din <= 32'h085ac6b6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ff; din <= 32'h87a6530e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h077; din <= 32'h8ff74e89;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h366; din <= 32'h1b1bacef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17c; din <= 32'h21e67dc7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1dd; din <= 32'h04a7abec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06f; din <= 32'he9c99763;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ec; din <= 32'hc8bed9df;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h373; din <= 32'hc12db33c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c9; din <= 32'h89953038;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h200; din <= 32'h7860ead0;

        // Finish
        @(posedge clk); en <= 0;  addr <= 10'hxxx; din <= 32'hxxxxxxxx;
        repeat (5) @(posedge clk);
        $finish();
    end

    always #1 clk = ~clk;
endmodule
