`timescale 1ns / 1ps

module testbench #(parameter DATA_WIDTH = 32, parameter BYTE_ADDR_WIDTH = 8, parameter BANKS_ADDR_WIDTH = 2);
    reg clk;
    reg en, wen;
    reg [BYTE_ADDR_WIDTH+BANKS_ADDR_WIDTH-1:0] addr;
    reg [DATA_WIDTH-1:0] din;
    wire [DATA_WIDTH-1:0] dout;

    seq_bank uut (
        .clk(clk),
        .en(en),
        .wen(wen),
        .addr(addr),
        .din(din),
        .dout(dout)
    );

    initial begin
        $dumpfile("waveform.vcd");
        // $dumpvars(0, testbench.uut.en, testbench.uut.wen, testbench.uut.addr, testbench.uut.din, testbench.uut.dout);
        $dumpvars(0, uut);

        // Initialize
        clk = 0;
        en = 0;
        wen = 0;
        @(posedge clk); en <= 0;
        @(posedge clk);

        // Autogenerated code        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d2; din <= 32'ha511ef01;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h038; din <= 32'h0eb328bb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e5; din <= 32'h1800d096;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07a; din <= 32'h166c05f1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15a; din <= 32'hf71b2096;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h057; din <= 32'h6d30bb2d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23b; din <= 32'he21b6fab;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h056; din <= 32'hcd088712;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32c; din <= 32'haae74af1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cd; din <= 32'ha1543af2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h191; din <= 32'h2a1f55b4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0af; din <= 32'ha3126780;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ff; din <= 32'h328ae691;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08d; din <= 32'h8fcf3c3f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h375; din <= 32'h713a702d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h098; din <= 32'h64f16362;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b9; din <= 32'ha63da8c8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h071; din <= 32'h3518a2e3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h232; din <= 32'h9ae1bdf3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h033; din <= 32'h724b7626;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34e; din <= 32'haeefa677;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09e; din <= 32'h09b580ce;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12d; din <= 32'he25d4004;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0aa; din <= 32'hbe8da94c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cb; din <= 32'habbd65d6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a4; din <= 32'h44fc11aa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37d; din <= 32'hb25ca15e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h096; din <= 32'hdfaf7c7b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h115; din <= 32'h68290d48;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09f; din <= 32'h0567f8da;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25b; din <= 32'he767cd28;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h086; din <= 32'h8b065783;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37b; din <= 32'hecc8252c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07c; din <= 32'h338adeb0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a0; din <= 32'h4f9d9a67;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a6; din <= 32'hb2f02895;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e3; din <= 32'h077597af;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h011; din <= 32'h7916a0a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fb; din <= 32'he77144ed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h067; din <= 32'h12ac9124;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h123; din <= 32'h43a0a487;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e8; din <= 32'hd1e7f2bd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f3; din <= 32'h0b0b8261;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h004; din <= 32'h058b0140;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3dc; din <= 32'h7a303f03;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h018; din <= 32'hde0dd98a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bc; din <= 32'habd378e2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h028; din <= 32'h2288d489;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24f; din <= 32'h37dbc198;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ac; din <= 32'h5ff0882a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b1; din <= 32'h8f0c8d23;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h069; din <= 32'h482e295c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18f; din <= 32'h5a7aa14a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h058; din <= 32'hb771bd99;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h247; din <= 32'h5931bdf3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d5; din <= 32'h4b7db429;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h396; din <= 32'h318af28d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h061; din <= 32'h8e1ca3bd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h130; din <= 32'ha464c414;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h037; din <= 32'h57112c17;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b9; din <= 32'h45380938;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ac; din <= 32'h04acfdc1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34f; din <= 32'hc250171f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b4; din <= 32'ha1c77a0f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13e; din <= 32'h771cb00b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h052; din <= 32'h8851e293;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h294; din <= 32'h850dfec1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04f; din <= 32'haaf445a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30c; din <= 32'h03e7a67a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10b; din <= 32'h61d24110;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c1; din <= 32'h53d05c70;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a6; din <= 32'h1f60aef8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h328; din <= 32'h7ff30bf0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17c; din <= 32'h73ef817a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h206; din <= 32'h4a0ffb46;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h096; din <= 32'hbf94743e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b3; din <= 32'h900a69b3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ad; din <= 32'h6f0382e6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f6; din <= 32'he24ae359;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03c; din <= 32'h4dd9f40a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ff; din <= 32'h547782c7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h183; din <= 32'hcb10c727;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h259; din <= 32'h5e666e59;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h054; din <= 32'h4693bafc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e6; din <= 32'h0d0a3efa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1df; din <= 32'h87eab583;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h234; din <= 32'h85bee34a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02b; din <= 32'h450c2352;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h386; din <= 32'h30cd7a43;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13b; din <= 32'hbfecb20a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h238; din <= 32'h8d83836d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h043; din <= 32'h3731e87a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3be; din <= 32'h75211d85;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h146; din <= 32'heb970d15;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h265; din <= 32'h92639b71;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h056; din <= 32'h6584f71a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c5; din <= 32'hf3b77501;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ea; din <= 32'h1643c058;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h273; din <= 32'h9196051b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h016; din <= 32'h4fb12ace;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f9; din <= 32'h7cbe2442;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h128; din <= 32'h715deee3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27e; din <= 32'hbdc200e7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d3; din <= 32'h933a4996;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f2; din <= 32'h04647eed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h114; din <= 32'h1bda904a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e0; din <= 32'hf9031555;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07c; din <= 32'hb4588a4a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ed; din <= 32'h54924618;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h138; din <= 32'hdb8a5eda;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ce; din <= 32'h580e2045;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fd; din <= 32'h7ad61d01;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ac; din <= 32'hf46ee485;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12f; din <= 32'h49f7eccf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2fe; din <= 32'h372da00b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0da; din <= 32'hd1fa9c3a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h373; din <= 32'h0d47843f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bd; din <= 32'h50f440e8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ca; din <= 32'h2ff27841;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h043; din <= 32'h6498abeb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h332; din <= 32'h616649b3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13c; din <= 32'hc35b1026;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h265; din <= 32'ha180a23a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c7; din <= 32'h7f10d4d4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h378; din <= 32'h034b8603;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13b; din <= 32'h3f8c5f37;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cd; din <= 32'hfc390461;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h082; din <= 32'h7b595c6a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h321; din <= 32'he3383e55;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h113; din <= 32'h4c139bbd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a4; din <= 32'h0d6db616;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02f; din <= 32'h975a3c5b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b3; din <= 32'ha319df6f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18d; din <= 32'h93500621;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h273; din <= 32'hd7f0829a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h043; din <= 32'h23361bfe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h377; din <= 32'h7cfc93e2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h185; din <= 32'h84904f53;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a4; din <= 32'h8adfca5e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08d; din <= 32'h71d995b9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h347; din <= 32'h4e772174;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16c; din <= 32'hee0f3ed0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28f; din <= 32'h3e6bc9e1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h013; din <= 32'h7bad80bd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e0; din <= 32'h54fe6670;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a7; din <= 32'he06985e3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22a; din <= 32'h2a2650a2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h072; din <= 32'h77ea101f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35e; din <= 32'h63df72aa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h177; din <= 32'h76c73c8c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h231; din <= 32'h02c6906f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04c; din <= 32'h31807f01;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h315; din <= 32'h09f767f3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h193; din <= 32'hfcfda714;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h275; din <= 32'h623a16eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e9; din <= 32'hdb24c403;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31a; din <= 32'h6e814153;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h150; din <= 32'hfaac46b3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20e; din <= 32'hb6b662b2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09a; din <= 32'ha9374b71;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34f; din <= 32'h33b8b48d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17f; din <= 32'h8e6f59c4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h291; din <= 32'h9229da34;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h019; din <= 32'h79c38e1b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h335; din <= 32'hd339d1d3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cc; din <= 32'h7ff29db5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h261; din <= 32'h2a13b842;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h077; din <= 32'h20fb030d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h359; din <= 32'h41e49732;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h143; din <= 32'h0641342c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h257; din <= 32'h33ebc5d6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d0; din <= 32'h6d77589a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h335; din <= 32'h260ff7d1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h160; din <= 32'hfdc88d56;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a6; din <= 32'hc15920fd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02f; din <= 32'he2457993;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d7; din <= 32'h92cdcc58;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h172; din <= 32'hc3d8c023;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h273; din <= 32'he73066af;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h095; din <= 32'he5b216f4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36a; din <= 32'h05db5d2d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ef; din <= 32'ha6556f58;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h201; din <= 32'hc7710f39;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fd; din <= 32'h763f64fc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h370; din <= 32'h73b721a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h119; din <= 32'hd445383f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h247; din <= 32'hccca434a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h018; din <= 32'h0966585e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h348; din <= 32'hcf578297;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16b; din <= 32'hf70a4ccc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24c; din <= 32'hcaf88877;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00e; din <= 32'ha55a468d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h336; din <= 32'h5cc73e66;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15c; din <= 32'hc63c8f6b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h235; din <= 32'hc99f34e1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05d; din <= 32'h623d2b54;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b0; din <= 32'hd9ac1c7f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h177; din <= 32'h2af2deaa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a4; din <= 32'h64da74d3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h091; din <= 32'hdc66b4e7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30c; din <= 32'h4cccd161;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h194; din <= 32'h5d1faae3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h230; din <= 32'h61df7f1b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h056; din <= 32'h6a93110a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34a; din <= 32'h1690c715;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h199; din <= 32'h5b752e9b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c5; din <= 32'hc1a1ff4e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05f; din <= 32'ha530eb3c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h327; din <= 32'h12b8464d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16c; din <= 32'h5329d2a8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e4; din <= 32'h94e5bb3c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03c; din <= 32'h5629cd4f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h393; din <= 32'h4a523b16;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18b; din <= 32'h06f7aaa4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b6; din <= 32'hb361423a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h045; din <= 32'h9e0ffd70;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38a; din <= 32'hf444ec2f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14f; din <= 32'h3af17cd9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ae; din <= 32'h71244423;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cb; din <= 32'ha86a2178;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a9; din <= 32'h0e75c70f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a7; din <= 32'h015e41d4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20e; din <= 32'h25fa3687;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h057; din <= 32'hef8c0074;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39f; din <= 32'h0aac4629;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ea; din <= 32'h70c4378b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h201; din <= 32'h7308d9d7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01f; din <= 32'hb4ade5cf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32a; din <= 32'hfb4b9051;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h159; din <= 32'h1d137251;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h247; din <= 32'he23d7fab;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ee; din <= 32'h81ad33fe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34c; din <= 32'hcf545f31;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h146; din <= 32'hbb5dd7af;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a6; din <= 32'h0cb1a994;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h027; din <= 32'hd92d97d4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33e; din <= 32'h178616b5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h133; din <= 32'h953868c5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h286; din <= 32'h1971ff47;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h056; din <= 32'h6b435b62;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a5; din <= 32'h321d7e05;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h163; din <= 32'h180d1051;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h250; din <= 32'h1271e93f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h061; din <= 32'h375894e7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h310; din <= 32'hff1548b4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h101; din <= 32'hd19fcf04;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a6; din <= 32'hd5bf6d4f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00f; din <= 32'hc298b762;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37c; din <= 32'h675d5b57;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ee; din <= 32'h019a7fe6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h220; din <= 32'h2b2414af;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a3; din <= 32'h1508935b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e1; din <= 32'h429b2671;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11a; din <= 32'h308a41a8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h262; din <= 32'hd9b75700;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h076; din <= 32'hc3b455ab;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37f; din <= 32'h337b1400;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f4; din <= 32'h79f87487;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bd; din <= 32'h6faae64e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d8; din <= 32'h392f8e5e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h301; din <= 32'h97d10c92;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h141; din <= 32'hedea24da;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ad; din <= 32'hd31ca524;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f6; din <= 32'hc8e6a67f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35b; din <= 32'h42366c2b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d0; din <= 32'hcb0204cc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cd; din <= 32'he008f6bd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bb; din <= 32'h55b36fd4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h320; din <= 32'he2414c08;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h164; din <= 32'hb16e7e92;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cd; din <= 32'h4d2b1a01;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04a; din <= 32'h0b4fd406;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h349; din <= 32'hf591d009;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h145; din <= 32'h6482b8e4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26d; din <= 32'h0ddf47fb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0aa; din <= 32'h39abd4fa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3de; din <= 32'hcd8012b7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h136; din <= 32'h63cb7060;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h291; din <= 32'h68332ffe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h056; din <= 32'hca0847a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h364; din <= 32'hd07144c6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15f; din <= 32'h7630f610;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h269; din <= 32'h924d0581;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h062; din <= 32'he2cfd409;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h318; din <= 32'h852c7426;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fc; din <= 32'h5486da98;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h251; din <= 32'h2afe9814;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02a; din <= 32'hd6d8ec47;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c6; din <= 32'hec206a02;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h132; din <= 32'hd04611b1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d8; din <= 32'h2684bd4d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h038; din <= 32'h22a71c15;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a3; din <= 32'hb6f57516;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h183; din <= 32'hede293bd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c5; din <= 32'hf66f8ead;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fd; din <= 32'h479d450b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ea; din <= 32'hcc9a7b07;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h133; din <= 32'h968d0b7d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h209; din <= 32'h2fe15a09;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08e; din <= 32'h9477403b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e8; din <= 32'ha0b7c34d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h176; din <= 32'hf2bc5db3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22c; din <= 32'h7ddec023;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c9; din <= 32'hd6b25be5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h350; din <= 32'h7b732663;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17a; din <= 32'hc09d8d93;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h228; din <= 32'h0ecf5112;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h032; din <= 32'h2afe964b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h332; din <= 32'h6cdb98b2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h171; din <= 32'h20b7621d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24a; din <= 32'h7e79f41e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e7; din <= 32'h0756001b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h395; din <= 32'h790c7aed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fd; din <= 32'ha5fe8a69;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h201; din <= 32'h612789c8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0af; din <= 32'h41d5a86e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h366; din <= 32'h4df011d1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d2; din <= 32'hdfe7dbc7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2fc; din <= 32'h2f9c8ed9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d9; din <= 32'h91b91104;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35e; din <= 32'he094fe93;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h114; din <= 32'hf40dc306;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26a; din <= 32'h15f11b05;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h065; din <= 32'hdca75a12;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d8; din <= 32'h0ad3c4cc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f3; din <= 32'ha657ecbd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ca; din <= 32'hb63d2d7e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09a; din <= 32'hfbbe05e0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h398; din <= 32'hff541025;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c7; din <= 32'hcab5fca2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23f; din <= 32'h5f037d02;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b4; din <= 32'hbba2dcb8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3df; din <= 32'hccbbbbb3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h152; din <= 32'ha77ccb61;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ce; din <= 32'h0edf831f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a8; din <= 32'hdcbb1037;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33d; din <= 32'h597c3da0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16c; din <= 32'h491575af;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24a; din <= 32'h9b56d76e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c7; din <= 32'hc25bb209;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34e; din <= 32'hd2176d9a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10d; din <= 32'ha6f132cd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h221; din <= 32'h13735318;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e9; din <= 32'hc1d8e770;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b6; din <= 32'h83c49ed2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c7; din <= 32'h438ed671;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h256; din <= 32'h102b4295;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h083; din <= 32'hfa6fa5fa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31f; din <= 32'he5785bb5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ef; din <= 32'h684a2863;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h205; din <= 32'ha5a2ffa3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04b; din <= 32'hdc5e1128;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32a; din <= 32'h039305f1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h118; din <= 32'h09a1bbab;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h247; din <= 32'h96108b2b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05d; din <= 32'he819eb25;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h363; din <= 32'h3563f25c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h150; din <= 32'h0a73c171;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22f; din <= 32'h2f643c33;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01d; din <= 32'h0c8e7137;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h346; din <= 32'h76cbfd69;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h100; din <= 32'h98780a2b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a2; din <= 32'h69fcad50;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h044; din <= 32'h20f8c87c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h344; din <= 32'hdb00d053;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h165; din <= 32'h1016383a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ce; din <= 32'ha21ee6ec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08c; din <= 32'hb681ed76;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e6; din <= 32'h9605116a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h138; din <= 32'h40c70f6d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cf; din <= 32'h0ed511c0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h016; din <= 32'hcb8a38c3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h358; din <= 32'h0e165c88;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11a; din <= 32'h7eb4519a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b4; din <= 32'h80b508eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b2; din <= 32'h18a6a96d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33e; din <= 32'he7148647;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c5; din <= 32'ha4b3a592;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e2; din <= 32'h86344a8f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ec; din <= 32'hd49320af;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31b; din <= 32'h9b2f4410;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18f; din <= 32'h59d9b69a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b5; din <= 32'hbe00e056;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f1; din <= 32'hf6fdfaae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h341; din <= 32'hb5ecbd8c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cc; din <= 32'hf87d5083;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2aa; din <= 32'h7201a079;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ee; din <= 32'hf47b0ee2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h388; din <= 32'h4327fbd7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18e; din <= 32'ha405510a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h252; din <= 32'h44e2cae2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bc; din <= 32'hce98faae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31b; din <= 32'h738d149c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18d; din <= 32'h5ec5cb9c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b9; din <= 32'hd17f3bf7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08a; din <= 32'h1d0719d2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3aa; din <= 32'h7c083df5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c0; din <= 32'h1b63eec9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ab; din <= 32'h4e294748;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02d; din <= 32'hf639c91f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h323; din <= 32'hd2a9d66f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1dc; din <= 32'h0e089d9d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h201; din <= 32'hdf16333e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a0; din <= 32'h2a4319f1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34c; din <= 32'hdea62b41;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b0; din <= 32'h52680ff8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h291; din <= 32'h6fe5989f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h020; din <= 32'h4fe1412c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36c; din <= 32'he028f645;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10e; din <= 32'h1153d83e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h253; din <= 32'h43f682dd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h056; din <= 32'hb98a391e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36e; din <= 32'h45cdf289;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h136; din <= 32'hb4fe12bc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h281; din <= 32'hd58709a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01e; din <= 32'h9c2240c8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h327; din <= 32'h31c294d8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h192; din <= 32'hd13c9fac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26d; din <= 32'hbc0385de;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03e; din <= 32'hb2957f01;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35e; din <= 32'h90297ef6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h115; din <= 32'h58bbef9a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h299; din <= 32'hf925a959;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06b; din <= 32'h5b304943;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e1; din <= 32'hb63a30ef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h119; din <= 32'hbc51b6d0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25f; din <= 32'hea82fc7b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b7; din <= 32'h834f235c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fe; din <= 32'h4dc65217;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h149; din <= 32'h928e31f0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h276; din <= 32'h51af9838;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01a; din <= 32'hae25a29a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35b; din <= 32'hc6655239;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ea; din <= 32'h65466e53;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h279; din <= 32'h9a282ac6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h088; din <= 32'h9ff52465;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d5; din <= 32'h6544d3f6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h137; din <= 32'h18162276;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h261; din <= 32'hf83e57b3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08e; din <= 32'haad8d5be;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35f; din <= 32'he2c4d782;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1df; din <= 32'h949cb614;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2fe; din <= 32'h7bd25426;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b3; din <= 32'ha2021a77;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e9; din <= 32'h604c4ed2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h101; din <= 32'hf54daff3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h204; din <= 32'h25a5e8f7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f7; din <= 32'h2ebb32f2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h316; din <= 32'h55f5d091;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bf; din <= 32'h69866baf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24a; din <= 32'h80dea921;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cb; din <= 32'h085622f5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39e; din <= 32'h4fcb7723;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d4; din <= 32'ha0573641;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2aa; din <= 32'h8062f1e6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cb; din <= 32'h68cf6b25;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h318; din <= 32'hc68c94c4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h150; din <= 32'hac66fc8b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2af; din <= 32'hddcb6620;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05d; din <= 32'h467434c7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c1; din <= 32'h09e346d5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19e; din <= 32'h34379642;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c4; din <= 32'h6f8551a5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03c; din <= 32'h0e17ddec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35a; din <= 32'h572b5e56;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1af; din <= 32'h83178309;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h282; din <= 32'h99c2b937;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h033; din <= 32'hd317cb1c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fb; din <= 32'h890e40c5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f0; din <= 32'h3e51c8aa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d0; din <= 32'hb0123e71;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h070; din <= 32'hb6b28986;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35f; din <= 32'heed1cbf6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18f; din <= 32'h2ae6a1a5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h277; din <= 32'h26043752;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ca; din <= 32'h931de439;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a7; din <= 32'h11b389af;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f9; din <= 32'hec64c9fa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f9; din <= 32'h29c40000;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09c; din <= 32'hecc1fffe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b1; din <= 32'h9b8ae312;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16f; din <= 32'h5e8a2cfe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2fe; din <= 32'h105eeb0e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07d; din <= 32'hba0623e1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ac; din <= 32'h5ad94432;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18d; din <= 32'h2fc6db26;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e2; din <= 32'hf585fe7d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h099; din <= 32'hd6940c91;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30e; din <= 32'h92928214;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h162; din <= 32'hcd0f6aeb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f4; din <= 32'h3a58a4b5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h037; din <= 32'hcce7eb3d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h394; din <= 32'h0fa051cb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h100; din <= 32'h61beb23e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22d; din <= 32'hc6ddc326;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h004; din <= 32'h62dd207a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37e; din <= 32'h8dc0bd29;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ef; din <= 32'h585359cc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f0; din <= 32'heecfc849;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01a; din <= 32'h33e3a588;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c4; din <= 32'hf845dae9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h178; din <= 32'he905a6d8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26e; din <= 32'h7017e5ee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h032; din <= 32'hc4a8a8b5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h311; din <= 32'he6fb16a9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ca; din <= 32'h7b5e6da1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24b; din <= 32'h33f12adf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h025; din <= 32'he017813d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h312; din <= 32'hd26e2c2b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15d; din <= 32'h2cb8af71;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c4; din <= 32'hfa56f363;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ac; din <= 32'h4b77b76f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3aa; din <= 32'h649a6913;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ce; din <= 32'h5c12cce0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h267; din <= 32'ha3040007;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h062; din <= 32'h84a01ca1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h327; din <= 32'h44210d44;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h104; din <= 32'h80ef18c5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e8; din <= 32'h2c56c653;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h060; din <= 32'h4ee3f352;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h397; din <= 32'hceed40a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17e; din <= 32'h67888581;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h245; din <= 32'h8b243883;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h027; din <= 32'h375b5da6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h372; din <= 32'h0582d76d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h174; din <= 32'h0c58115f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h263; din <= 32'hf53ffd64;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b8; din <= 32'h9afc25e7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39a; din <= 32'hfd1449f0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h101; din <= 32'h0299091e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h234; din <= 32'hff135121;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h096; din <= 32'h0c343f67;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39f; din <= 32'h4526e5b4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e2; din <= 32'hfbadb724;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h225; din <= 32'hbdefbeeb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08c; din <= 32'h124049e1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f7; din <= 32'hf52b937e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1be; din <= 32'hae62f44e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c4; din <= 32'hb92d4c9b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d8; din <= 32'hf07998dc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ba; din <= 32'hf8b37304;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h131; din <= 32'hbc4d5c66;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25f; din <= 32'hc4f2b84b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0aa; din <= 32'h41665bae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ed; din <= 32'hf67e07f9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12e; din <= 32'h8e946cea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21b; din <= 32'hf32d40cb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07f; din <= 32'h554d2c5a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3eb; din <= 32'h57aa6bd8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h148; din <= 32'h4cc91f6c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h274; din <= 32'h29c9ad1b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c3; din <= 32'hde92a080;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h314; din <= 32'hc7ea0717;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h163; din <= 32'h39f7fbdc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h209; din <= 32'hd21c4a7c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ac; din <= 32'h962ec1df;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h382; din <= 32'h342bbf77;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h113; din <= 32'h3a701330;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h257; din <= 32'hc2ac0b27;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a2; din <= 32'he4732e94;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30b; din <= 32'hfc3e219c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h129; din <= 32'h6d70a845;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29a; din <= 32'h4c525a5f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h079; din <= 32'hf6bcf122;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35f; din <= 32'h952e4356;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f3; din <= 32'h50501e90;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20e; din <= 32'h4f2be303;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a2; din <= 32'h45baa30c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fc; din <= 32'hf3d9c3d3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a6; din <= 32'h11c596dd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23e; din <= 32'hbb6103b5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h046; din <= 32'h1a81fcc3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h322; din <= 32'hc81f7651;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bd; din <= 32'hdf76bcd5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h241; din <= 32'h33141ed1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b7; din <= 32'h47438082;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39d; din <= 32'h9643c50c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h113; din <= 32'h9534cc3c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h214; din <= 32'h434ef346;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h069; din <= 32'hc1373ecd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h338; din <= 32'h854b47c8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1de; din <= 32'h4bf6dbd2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ed; din <= 32'h2ef4c45a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f6; din <= 32'h8f619bf9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h358; din <= 32'h7d80b42d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11e; din <= 32'hff9d07a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h290; din <= 32'hc5cf0848;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b3; din <= 32'ha20ca5f8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30f; din <= 32'hb1e7d9a2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h186; din <= 32'h5bb44395;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ab; din <= 32'h6ef175ec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0de; din <= 32'h1f86d44c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32f; din <= 32'h8c2bb188;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1aa; din <= 32'hc3c0ef20;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e9; din <= 32'hd69079b6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09e; din <= 32'h4fdae04d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h390; din <= 32'h1c7ee31e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11b; din <= 32'hf190d15c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h259; din <= 32'h1697ef88;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08f; din <= 32'hba32253b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h320; din <= 32'ha2bbf170;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18d; din <= 32'h1c56a3f2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h292; din <= 32'h68e01a3f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bc; din <= 32'h82e2909b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30b; din <= 32'h3cebd937;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h118; din <= 32'h6ee45df5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23f; din <= 32'h7e6f7123;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h045; din <= 32'hd61cfb06;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34f; din <= 32'h8c21fd39;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h110; din <= 32'hf5a5086d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22a; din <= 32'h21a86fe9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h081; din <= 32'hf8f80777;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a2; din <= 32'h3b264eb2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h188; din <= 32'h18eae9a4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bb; din <= 32'ha79b4ff4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09a; din <= 32'h284b71ce;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h325; din <= 32'h3d3a8adf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d7; din <= 32'h425f7f22;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h201; din <= 32'h2592478d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00c; din <= 32'hb8782294;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36b; din <= 32'h3731fdaf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d0; din <= 32'h2f52185b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2db; din <= 32'h89d65146;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h048; din <= 32'h788eae8c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f1; din <= 32'h5900e5a1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e3; din <= 32'h86e8e6f0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h264; din <= 32'h0b91182c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h037; din <= 32'hf8fecae1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h309; din <= 32'h85cfb50b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h132; din <= 32'h4c4a3bd4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22f; din <= 32'h91eb8324;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h003; din <= 32'h9d875818;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c7; din <= 32'hd1c702a7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h180; din <= 32'h46f10883;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b6; din <= 32'h0f3f0995;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ec; din <= 32'hc1ded558;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d5; din <= 32'hd8f55b1b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h135; din <= 32'hae2e7ebd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c5; din <= 32'hf1fc3fd9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cc; din <= 32'h176196d0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ca; din <= 32'h26c073be;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a5; din <= 32'hf6f96aba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h290; din <= 32'hb9491b06;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h072; din <= 32'h58fc546e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36b; din <= 32'hec10704b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f4; din <= 32'h3dab8c0d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ca; din <= 32'h3489d82f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00d; din <= 32'h5fd23a87;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h301; din <= 32'h6ea8cf40;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15e; din <= 32'h3009953c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ee; din <= 32'he2d0bc6c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e0; din <= 32'h56ce2229;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35d; din <= 32'h1c43ee1b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13b; din <= 32'h5bdda68d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h215; din <= 32'h68634ffd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h077; din <= 32'hcb0a196c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h354; din <= 32'h2c826741;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h169; din <= 32'h0ebdf3b6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h220; din <= 32'he9b8d548;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e4; din <= 32'haa89295f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h325; din <= 32'hd07adbfe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10a; din <= 32'hd77bb47f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26b; din <= 32'h1fafe22e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fd; din <= 32'h702ebbc3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d7; din <= 32'hf86fe731;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h180; din <= 32'h22f1c370;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cf; din <= 32'hc56fc99c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06a; din <= 32'hb6746025;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ad; din <= 32'ha5108bc8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h179; din <= 32'he6ee45dc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h285; din <= 32'h10e4bb17;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h043; din <= 32'h97b56aa7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33e; din <= 32'hd7cd9c54;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h115; din <= 32'hb65e387b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ab; din <= 32'hef77d9d9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b2; din <= 32'hd960a690;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37d; din <= 32'hf28d013e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e5; din <= 32'h0f230895;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h291; din <= 32'hfecdcfea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0dc; din <= 32'h89179fd2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39f; din <= 32'hc004388a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11d; din <= 32'h53e1402b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2da; din <= 32'h651ee498;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h027; din <= 32'he15ed7a5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33b; din <= 32'h65cdd0c1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d9; din <= 32'h02ed5ded;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20f; din <= 32'he8859a07;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06c; din <= 32'hb67e1efa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h342; din <= 32'h38fb995d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12e; din <= 32'h28108eeb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21f; din <= 32'h3dcf10ca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d8; din <= 32'h97fb060f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e2; din <= 32'hace01afe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fe; din <= 32'h690cdbab;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b0; din <= 32'hb9b6e30b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c2; din <= 32'h930bc5c0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h309; din <= 32'h512d0382;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h121; din <= 32'habd1c579;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2db; din <= 32'hdd485db6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d5; din <= 32'hf4ee01cf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h327; din <= 32'h1873b6ea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h170; din <= 32'h2b047b5a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f4; din <= 32'h168c5683;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0eb; din <= 32'h211eae88;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h390; din <= 32'hcf530a1a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a8; din <= 32'h24359580;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23e; din <= 32'h40c92798;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00b; din <= 32'h28181f1e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e0; din <= 32'h45582322;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fe; din <= 32'h0fecb1a5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a8; din <= 32'hd697b4e2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h018; din <= 32'h21e3e673;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h337; din <= 32'h84b35ec6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h164; din <= 32'hb207729d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a2; din <= 32'h6505cc7b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h089; din <= 32'h4b9948e3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h314; din <= 32'hf0e0c71f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12c; din <= 32'h34eea130;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a5; din <= 32'h2a928f16;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0de; din <= 32'h0b03a7a1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39b; din <= 32'h0e608121;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10c; din <= 32'hd6f2e758;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h297; din <= 32'h957c6a06;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08d; din <= 32'h82181338;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d7; din <= 32'hdce9fd8a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19f; din <= 32'hff7c1b37;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b3; din <= 32'hb3fb62b8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a6; din <= 32'h77ab688f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ac; din <= 32'hb2c1a35a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h160; din <= 32'h31924001;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h231; din <= 32'hb3a947c3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05e; din <= 32'ha7b65810;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h365; din <= 32'h0983123f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h162; din <= 32'hc7fcd1aa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22d; din <= 32'hc60c1d4f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ac; din <= 32'h95ba5503;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h362; din <= 32'h8cb69c36;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1af; din <= 32'h21922628;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26f; din <= 32'h492865f5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h065; din <= 32'h00ee1e05;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35e; din <= 32'hf8873b50;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h163; din <= 32'h64fc9f1d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27f; din <= 32'haa9779d6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fe; din <= 32'hc925c52e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h308; din <= 32'hab4a680d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15e; din <= 32'hd703804e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22d; din <= 32'hb55bf8ab;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d0; din <= 32'hd3fdc1ff;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d9; din <= 32'h7e704315;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h186; din <= 32'hecfa2884;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h219; din <= 32'h59766461;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a3; din <= 32'hfb5763cb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h371; din <= 32'h53738342;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h134; din <= 32'h1d4fcc89;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2df; din <= 32'he462f5b0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h092; din <= 32'hf02ccffc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h365; din <= 32'hf01ddfea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b3; din <= 32'h7fee228b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22a; din <= 32'h72c0f9f3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e7; din <= 32'h797eff2f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h318; din <= 32'hd9226e70;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h199; din <= 32'h6e26e65a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27b; din <= 32'h6688335d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h049; din <= 32'h0f8c425c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f6; din <= 32'h5cf57011;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f0; din <= 32'h32125c46;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h266; din <= 32'h81c0f531;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h045; din <= 32'ha7b80794;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f8; din <= 32'h55bafcd2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16a; din <= 32'h0bfd850c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e3; din <= 32'hc91af1d6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b0; din <= 32'h371c580c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h357; din <= 32'hb9370f1b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c1; din <= 32'h4f149e83;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h231; din <= 32'ha9c3937a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cc; din <= 32'hbf4134dc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e4; din <= 32'he6e0a876;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1df; din <= 32'h1b111102;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a4; din <= 32'h070a7cc7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h010; din <= 32'h21b7257a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39a; din <= 32'h07185d04;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h140; din <= 32'h21b93647;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h256; din <= 32'h4c6e6686;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08a; din <= 32'h4aade046;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h315; din <= 32'habba810a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10c; din <= 32'h925a3a6f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h286; din <= 32'h53ff601f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ac; din <= 32'h70bdf19e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h366; din <= 32'h7a4c1c47;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h130; din <= 32'h57899f58;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cb; din <= 32'hc81ff5a7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a7; din <= 32'h0ad6abc4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h312; din <= 32'hb860b9b5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f3; din <= 32'h556fa401;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h212; din <= 32'h0e92fcd9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f9; din <= 32'ha6448b2c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e7; din <= 32'h5ae90231;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14d; din <= 32'h0e3579c3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26f; din <= 32'h6f8f695e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ec; din <= 32'h4398a392;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e2; din <= 32'h09a5ecaf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h188; din <= 32'hc728dd45;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h294; din <= 32'hd934b1ab;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e5; din <= 32'h12e561d3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b3; din <= 32'hb66bee94;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ed; din <= 32'h04f1f96d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ae; din <= 32'h8399769b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a6; din <= 32'he9452a71;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h368; din <= 32'h95264e80;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h129; din <= 32'hfd2ecd7b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20e; din <= 32'ha3d1e52d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a5; din <= 32'h7a7960ef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h361; din <= 32'h25cd2111;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h108; din <= 32'h81b65bd7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d6; din <= 32'hf2c5128b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h090; din <= 32'hab9fb9ed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h367; din <= 32'h3e28950b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h103; din <= 32'h861481cd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h241; din <= 32'h0640cdf8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h009; din <= 32'hd865a766;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h374; din <= 32'h7edf9c4c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a0; din <= 32'hafb4f8ad;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h295; din <= 32'hbb514264;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00d; din <= 32'hdc605a2a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h336; din <= 32'hd41b4774;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e3; din <= 32'h651b19b1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21c; din <= 32'ha9ddad82;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h089; din <= 32'h393c83a7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f2; din <= 32'h2985f6ba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h118; din <= 32'h8efd69c2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h287; din <= 32'h120c13e1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h063; din <= 32'h85b68fbe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h397; din <= 32'had3d8b02;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h192; din <= 32'hba033bca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b5; din <= 32'hab65b9eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b5; din <= 32'h99d660cd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b8; din <= 32'h4c85cb2c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d5; din <= 32'h2b384375;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f7; din <= 32'h4cb60df3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h095; din <= 32'h1073d107;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h366; din <= 32'h65ed3dd9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e3; din <= 32'h7223cebf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h259; din <= 32'h24ab46a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0de; din <= 32'h7c756772;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h304; din <= 32'h101f350b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h145; din <= 32'h14149a29;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h212; din <= 32'ha01800a8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d5; din <= 32'haa0c122e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b5; din <= 32'had4e2f67;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h141; din <= 32'ha80c55a8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25d; din <= 32'h9dbbd5f5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f0; din <= 32'hfebeb4f8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cb; din <= 32'h8fbf10dd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h126; din <= 32'hadf41f7e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a7; din <= 32'h7e446a6a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h023; din <= 32'h99c665b8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h320; din <= 32'hdab3d398;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d4; din <= 32'h98adce10;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cc; din <= 32'hd0e4f80d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ba; din <= 32'h3674b364;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33a; din <= 32'h3d60fd67;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h186; din <= 32'h2e48e1a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f4; din <= 32'hff8bec89;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h037; din <= 32'h297ad9f3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39f; din <= 32'habd1586a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d6; din <= 32'h0da93bf8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h282; din <= 32'h086ec43b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ab; din <= 32'hea1813bc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h394; din <= 32'hfe180f38;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h119; din <= 32'h56bb211a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h254; din <= 32'hfa7779f5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h072; din <= 32'h5a0884ff;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h380; din <= 32'hbab593ae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14d; din <= 32'hfd53d569;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h277; din <= 32'hf5c30680;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h049; din <= 32'hbd89af95;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h317; din <= 32'hed2d02b9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h183; din <= 32'h7f8ca5a7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d8; din <= 32'hdfb9f768;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06b; din <= 32'hd5118def;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h372; din <= 32'hcb715843;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14a; din <= 32'ha8a551eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h220; din <= 32'h74e6d48f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h016; din <= 32'ha92afa5d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32e; din <= 32'h6a9f35de;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h170; din <= 32'h0de101c8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2fe; din <= 32'hf32b4ee5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04d; din <= 32'hf61e63ba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d4; din <= 32'h9495bf02;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12a; din <= 32'h0dad27a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h218; din <= 32'ha2ee9438;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09c; din <= 32'h1cfef95e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39b; din <= 32'h464fce5e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12e; din <= 32'headae7e2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h286; din <= 32'h64a5f24e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h047; din <= 32'h7d9e39a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bd; din <= 32'hf03b1a85;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h113; din <= 32'h3ee0aaf6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e2; din <= 32'he59dffbb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00c; din <= 32'h147b6f07;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f6; din <= 32'h6ee65739;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h152; din <= 32'ha670be5e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e6; din <= 32'h6882ae49;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h007; din <= 32'h3ae57de8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h387; din <= 32'hcfd54150;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h117; din <= 32'hafff7f8b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26a; din <= 32'h23c3f8a7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h001; din <= 32'h690816f1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c1; din <= 32'hc33f334a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h102; din <= 32'h12f71436;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h238; din <= 32'hddbdee5c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h014; din <= 32'h22fe3dd4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e6; din <= 32'h15252aac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fe; din <= 32'h507938cb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22c; din <= 32'h3357520e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09e; din <= 32'hfcb38c19;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h397; din <= 32'h09e6d93e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a8; din <= 32'hfcddb024;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21c; din <= 32'h4af50f0e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09d; din <= 32'h1db91759;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ff; din <= 32'h456243cb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d9; din <= 32'hff267da6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23f; din <= 32'hcdafff5d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h087; din <= 32'h96419079;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e4; din <= 32'h20006fba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ab; din <= 32'h851bb3a8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h266; din <= 32'h290bd318;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h061; din <= 32'h040e8825;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d9; din <= 32'haa29c036;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c9; din <= 32'h1270931a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h234; din <= 32'hc5e0dfd5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ba; din <= 32'h488bb394;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h327; din <= 32'h9b77bfdc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18b; din <= 32'hc06d9f39;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d7; din <= 32'h35163e40;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h084; din <= 32'hb439fdc7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h301; din <= 32'h97f17841;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h174; din <= 32'hcfe80ab6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23f; din <= 32'hfb371325;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h000; din <= 32'hf7816fc6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h373; din <= 32'hadbf5fe3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h168; din <= 32'h60b6a595;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cf; din <= 32'h024d3548;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h090; din <= 32'hb99164e4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h365; din <= 32'h1a17964a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b7; din <= 32'he48b49f0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29d; din <= 32'h32878526;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c9; din <= 32'h121cf489;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f4; din <= 32'h073c8ebb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bb; din <= 32'ha649e5d6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d6; din <= 32'hdc1d8c59;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03c; din <= 32'h5b7fbd26;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h395; din <= 32'h05f825ec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cf; din <= 32'ha97af3f6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h252; din <= 32'hbc6c3092;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h065; din <= 32'h5162c23e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h383; din <= 32'h45251eab;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h109; din <= 32'h7d0cefb8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ea; din <= 32'hd95319ef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ce; din <= 32'h4a1df12a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31f; din <= 32'h46b6ba19;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h116; din <= 32'h89473582;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28a; din <= 32'ha5aaad4b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a9; din <= 32'h55ad82f3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h372; din <= 32'h547e82da;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e3; din <= 32'hcd3ed88e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23b; din <= 32'h1adc5e9c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a4; din <= 32'hfdf4eebe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b5; din <= 32'h3bfb2b87;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a8; din <= 32'h88c8fadb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h280; din <= 32'h1f60d988;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h078; din <= 32'h1a38e7c9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h391; din <= 32'h5fb04f77;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h179; din <= 32'ha82cb2bf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ae; din <= 32'h0a52890c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h092; din <= 32'h935d7dd7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h380; din <= 32'h91d654a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f2; din <= 32'hec2a813b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h252; din <= 32'h1b4d851a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h061; din <= 32'h0450396e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39e; din <= 32'he22244a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h153; din <= 32'h8986945d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a4; din <= 32'h74dcbe24;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h042; din <= 32'h43529667;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b7; din <= 32'h0a57be7b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17c; din <= 32'h2a3906e7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h217; din <= 32'h5ce21f76;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h000; din <= 32'h02b60cce;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h310; din <= 32'h1c6a6c30;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d5; din <= 32'h36a7c5a3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b6; din <= 32'hc8a6a3c7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01f; din <= 32'h4d09da78;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d9; din <= 32'h6db5dbc5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e9; din <= 32'hc7a4de12;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h241; din <= 32'h791493db;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04d; din <= 32'h9b66d772;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37f; din <= 32'hadee445d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d2; din <= 32'haeae836b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23b; din <= 32'h75bf6c25;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0db; din <= 32'hfa59df2e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h398; din <= 32'hc922dfb4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h126; din <= 32'h6bf141e3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c7; din <= 32'h29d52424;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h076; din <= 32'hafd2fabb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32e; din <= 32'hb05bdfb9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h122; din <= 32'h06da8803;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ce; din <= 32'h75b30fd7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e6; din <= 32'h0a57dd58;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e3; din <= 32'h25d98dbe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d2; din <= 32'h79e630f5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f5; din <= 32'h2ab54486;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h063; din <= 32'h7e1f332b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3df; din <= 32'ha4430279;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f5; din <= 32'he6d3cc33;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f6; din <= 32'h5ee40daf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c7; din <= 32'he04a2420;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e2; din <= 32'h3f03735a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13a; din <= 32'h032da4ad;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c7; din <= 32'h8eba0f33;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d6; din <= 32'hc1a342a9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3dd; din <= 32'h187c4a84;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h193; din <= 32'h1d9a40c7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h269; din <= 32'ha74ec141;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cc; din <= 32'h3cd4a131;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32b; din <= 32'h5fc8a885;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h136; din <= 32'hcb82be19;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ac; din <= 32'ha348f09e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h051; din <= 32'heb28140e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h339; din <= 32'h9c568ed9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h102; din <= 32'h3fa89619;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d8; din <= 32'h3f244d20;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h014; din <= 32'h63ad0ced;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h358; din <= 32'h594d7f55;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1aa; din <= 32'h6b339490;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h218; din <= 32'h97a17255;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h047; din <= 32'h8f9f7324;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bf; din <= 32'h9eb9b22a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h147; din <= 32'hc02890e4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27d; din <= 32'h83e2edb2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02a; din <= 32'h909059e7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30a; din <= 32'haaa0bec4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h163; din <= 32'h5bea4417;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c0; din <= 32'h6d169909;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h058; din <= 32'h85fbf982;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38c; din <= 32'hbe83ab4a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h199; din <= 32'h3722ec30;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c5; din <= 32'h27ce28eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h043; din <= 32'h45bf5250;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a0; din <= 32'hedeb4712;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11d; din <= 32'h00436089;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29e; din <= 32'h9193adfb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04c; din <= 32'hb9ca8969;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ba; din <= 32'hd4a67270;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1dc; din <= 32'h79bbffc6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a8; din <= 32'h6a5a7056;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b4; din <= 32'h517bad9e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e6; din <= 32'hc2053f13;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h109; din <= 32'ha228cb94;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22d; din <= 32'h8fdaf97f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h027; din <= 32'hdb3b0f19;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c9; din <= 32'hb02323b1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h120; din <= 32'hc39fe688;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c7; din <= 32'h528758c2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04d; din <= 32'hae5114ed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b3; din <= 32'h9640d355;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f7; din <= 32'he15337b4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2dd; din <= 32'h7b3623a2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cb; din <= 32'hbef70952;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32b; din <= 32'h7aa2c49d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18a; din <= 32'h52d59caf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h288; din <= 32'hd4c5c597;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c6; din <= 32'hbda1696e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h359; din <= 32'h07d8370b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h171; din <= 32'h960220bd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24b; din <= 32'h5d50d059;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h019; din <= 32'h052db02e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bd; din <= 32'h7f79921d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h137; din <= 32'hf9770839;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28f; din <= 32'h6c120dc0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f2; din <= 32'h6243d3f4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b2; din <= 32'h3d2a90dc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f1; din <= 32'h1c9c381a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28d; din <= 32'h5891cf10;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09c; din <= 32'h20259adf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h300; din <= 32'h16407508;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h145; din <= 32'h46057249;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2dc; din <= 32'h218d1e75;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h069; din <= 32'he844b5cc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f9; din <= 32'h27ed3c79;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cd; din <= 32'h71b45bae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d4; din <= 32'h385c4638;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e1; din <= 32'h9d9ef9b5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h359; din <= 32'hb9803700;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h165; din <= 32'h681339d5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h294; din <= 32'hed08eec6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c0; din <= 32'hb208a002;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h324; din <= 32'hf2e9f57d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c6; din <= 32'h24015ee2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h220; din <= 32'h39c259d3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a0; din <= 32'ha0b86852;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h301; din <= 32'he9eea442;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h157; din <= 32'hb1552499;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e1; din <= 32'h74c032e8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h013; din <= 32'h62eb9d32;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b4; din <= 32'hf65c0729;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b4; din <= 32'h08325410;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h231; din <= 32'h18cf3046;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e9; din <= 32'h8c294e5e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e0; din <= 32'h6f5150bf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d9; din <= 32'h784155a5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2af; din <= 32'h434c2480;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02f; din <= 32'h88534449;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h336; din <= 32'heae7b0ee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16b; din <= 32'h74c5dcac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h292; din <= 32'h1162bbd6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e1; din <= 32'h3dd9d3d7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36a; din <= 32'h3de0cc2a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h138; din <= 32'h5aae4df5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d5; din <= 32'hfda77f2e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05f; din <= 32'h0bcd667a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d6; din <= 32'h63d20721;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h165; din <= 32'hca96ea7d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23e; din <= 32'h962998bb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h004; din <= 32'hd14b393f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d5; din <= 32'h834b9618;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18a; din <= 32'h88c3d1c2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h207; din <= 32'h4b0c350e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h042; din <= 32'h97643593;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h340; din <= 32'h420ff785;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h103; din <= 32'h81c56b40;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20b; din <= 32'h13e51241;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h067; din <= 32'h849ce86a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a1; din <= 32'h29ef0698;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b9; din <= 32'h837ad8b9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d0; din <= 32'hbc307d48;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0eb; din <= 32'h1c571917;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h302; din <= 32'hdf136e69;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14b; din <= 32'h79a38c18;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h258; din <= 32'hac03db64;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e4; din <= 32'hb817a42d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c8; din <= 32'hc97a83ac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h196; din <= 32'hccc7cf33;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22f; din <= 32'hcce0da04;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cc; din <= 32'hd0043b31;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37b; din <= 32'hb9bb695f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h139; din <= 32'he74de598;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a7; din <= 32'hcc6e54f7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e0; din <= 32'h0b91583c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e4; din <= 32'h042f699b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d9; din <= 32'hf0946153;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h266; din <= 32'hbd23d745;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h090; din <= 32'hb0e3a621;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32f; din <= 32'h51bad099;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h158; din <= 32'h06401694;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h218; din <= 32'h32c1dfac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h088; din <= 32'h183d5899;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34b; din <= 32'h562da6c9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12d; din <= 32'h68e168e8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b0; din <= 32'h25c8fa84;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ec; din <= 32'h77367f42;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h382; din <= 32'h5baa5a6f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h198; din <= 32'h222db0ca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20f; din <= 32'h5e5c51a8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ea; din <= 32'hc91edf9d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36b; din <= 32'h4d9559d0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h150; din <= 32'h4037d46c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e9; din <= 32'hbb7fcfe6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h057; din <= 32'h065a282f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34b; din <= 32'h67b27ee9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h101; din <= 32'hba185276;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h204; din <= 32'hc7735842;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06c; din <= 32'h2af5aba0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33f; din <= 32'hae42233d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b7; din <= 32'h03d6bbb2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c3; din <= 32'h3a770885;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09d; din <= 32'hf5ce7d54;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h302; din <= 32'hae054c08;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c7; din <= 32'h31e8c6cd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e0; din <= 32'hef91e7a5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07f; din <= 32'hda43a496;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32d; din <= 32'h2a88ac2e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d9; din <= 32'h93686a71;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23a; din <= 32'h55c28be9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d3; din <= 32'hc1e51229;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h369; din <= 32'hace0a397;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h138; din <= 32'h0f82f0ba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e5; din <= 32'h2ec66d35;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f7; din <= 32'h11d5fe3e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h308; din <= 32'hcbb107ae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b3; din <= 32'hee9087ef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26a; din <= 32'hb50150b2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f0; din <= 32'h40d3b313;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31a; din <= 32'hf5a6c0c9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h126; din <= 32'h88435550;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h240; din <= 32'h4a59f244;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09c; din <= 32'hc53e755e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e9; din <= 32'hd5100b14;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h130; din <= 32'hcc74b066;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26e; din <= 32'h232e28c9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h048; din <= 32'hab7b1498;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f9; din <= 32'h1864836a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h195; din <= 32'h100b6479;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ca; din <= 32'h18df157e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b9; din <= 32'h1f05df5e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37b; din <= 32'hec1e0abb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ff; din <= 32'h83795809;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20e; din <= 32'h9687639a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f3; din <= 32'ha648f446;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32f; din <= 32'h864e803c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19f; din <= 32'h8bfccd75;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b6; din <= 32'h75ec6904;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0aa; din <= 32'h6fd4f6c8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37b; din <= 32'h269b4eaa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15b; din <= 32'hab4ea6c4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h217; din <= 32'h36882650;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fa; din <= 32'he0783b08;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3dd; din <= 32'h029f2357;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d6; din <= 32'ha1d8f3c3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d9; din <= 32'h8fb75c81;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07d; din <= 32'hd4ad3d59;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38e; din <= 32'h199a2424;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19e; din <= 32'hf4ee76ea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bc; din <= 32'h52cfae4a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h030; din <= 32'hb0b32bbf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h303; din <= 32'h48305a04;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fe; din <= 32'h91a9caaa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28c; din <= 32'hcfb03572;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c2; din <= 32'h9809b092;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36f; din <= 32'h3ecf029c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h184; din <= 32'h08c01970;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h224; din <= 32'h5a89e879;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0aa; din <= 32'h99790e12;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a4; din <= 32'h2116509f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c2; din <= 32'h1f348f3c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h281; din <= 32'h08e869d4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h031; din <= 32'h1a14d785;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h336; din <= 32'hd0386fdc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h153; din <= 32'ha1e98a3f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f1; din <= 32'h207d332d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h082; din <= 32'hd882a927;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h344; din <= 32'h09189374;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h163; din <= 32'hc334bc17;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h255; din <= 32'h7faf339f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h045; din <= 32'h98e5aff9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h375; din <= 32'h188acde8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b8; din <= 32'h5a425cd3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22c; din <= 32'hb38ac35c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ac; din <= 32'h764c9e47;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36d; din <= 32'h27b05b8e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h177; din <= 32'hf1807c7f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cf; din <= 32'h3ecf09ca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f3; din <= 32'h27062fa1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h344; din <= 32'hcdbce2d8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19d; din <= 32'ha0e2d56e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h286; din <= 32'h7e3cf2bb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05d; din <= 32'h0ef056ca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h330; din <= 32'hc0eb4bfc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d0; din <= 32'ha6007752;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21f; din <= 32'h0b25e9b0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02c; din <= 32'h0b8ddbd6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h371; din <= 32'h9067aff9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11d; din <= 32'h563ca7c0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h291; din <= 32'haee7bb64;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f9; din <= 32'h2daf8ecf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ff; din <= 32'hfd61d0fc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fa; din <= 32'h3d2ea5e6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h244; din <= 32'h87fa4c04;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ec; din <= 32'h87300f76;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h384; din <= 32'h1e82da1e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fe; din <= 32'h8dc4040f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27d; din <= 32'hf6232604;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03e; din <= 32'h8382a83c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d3; din <= 32'hb91ebe86;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c3; din <= 32'h48fb2772;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h270; din <= 32'h91f4456c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h009; din <= 32'h069ae906;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bf; din <= 32'h46c94b73;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h140; din <= 32'h694f31aa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h295; din <= 32'h3a6ff3e4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h071; din <= 32'h9900abc9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h362; din <= 32'ha8fb191a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bb; din <= 32'hd37a43cd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h257; din <= 32'h9032ac7d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h014; din <= 32'hebe55b23;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36e; din <= 32'h0200fb78;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d6; din <= 32'h60b38b67;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c3; din <= 32'hff4b6a45;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04e; din <= 32'h06568662;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d8; din <= 32'h04a52f77;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14e; din <= 32'h24e1f9d5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27d; din <= 32'h70715774;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cd; din <= 32'hdd31dc06;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38b; din <= 32'hac530e4e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c7; din <= 32'hadada3e3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ad; din <= 32'h5b425828;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h083; din <= 32'hd4532dd4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35f; din <= 32'ha3d18aba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cd; din <= 32'h19f60ff9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27a; din <= 32'hdc61156b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h065; din <= 32'ha373990e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h321; din <= 32'h5a0dd21f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h151; din <= 32'h4a48e46b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21c; din <= 32'h9767f98b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cd; din <= 32'ha6d63a85;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h346; din <= 32'h2c524784;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h153; din <= 32'ha17b93c6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24b; din <= 32'h290d2c86;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h005; din <= 32'hba98e17f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h389; din <= 32'h38477308;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h170; din <= 32'h12c05e49;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h270; din <= 32'h9785f806;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ba; din <= 32'h2d58f9aa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h302; din <= 32'h3fc203fe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a8; din <= 32'hb2ca6336;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h219; din <= 32'h0517b2bf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h017; din <= 32'h29876c14;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a8; din <= 32'h7bd558a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h121; din <= 32'hd831d378;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27b; din <= 32'hb0528d5c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0dc; din <= 32'h76c69cf6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c3; din <= 32'h5f091430;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c5; din <= 32'h375d4c12;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h241; din <= 32'h1e89833f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h097; din <= 32'h7fde0fb4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34e; din <= 32'h337e8b5d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b1; din <= 32'h7912eb4a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bf; din <= 32'hf6f0854c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h097; din <= 32'hb40cb1a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3aa; din <= 32'hd7e611c1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h104; din <= 32'h6727b401;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24f; din <= 32'hd845dec3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b4; din <= 32'hf273b8e3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39a; din <= 32'h36522ee4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h184; din <= 32'h98d70e80;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h239; din <= 32'heacd7407;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h084; din <= 32'h5d96dcfe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h327; din <= 32'hedf3ec7a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1aa; din <= 32'h5c729a7d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e0; din <= 32'h0cab1a6c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h092; din <= 32'hf21a3134;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h372; din <= 32'h67e32615;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h107; din <= 32'he392a12e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b0; din <= 32'hde4103de;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h059; din <= 32'hd2b22b55;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37d; din <= 32'hbb0c92c7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h132; din <= 32'hb1cce428;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22e; din <= 32'hfe08bcfe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07c; din <= 32'ha26e68fc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h388; din <= 32'ha5c565ad;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ab; din <= 32'h42c2c33b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h297; din <= 32'hbefd47b8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0da; din <= 32'hd8721497;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h306; din <= 32'h92674c90;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h129; din <= 32'hf7da02cc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bd; din <= 32'haa5e7300;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05c; din <= 32'h91ea134e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33d; din <= 32'h092462b0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h125; din <= 32'h68a65102;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h201; din <= 32'h41ca2edf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a2; din <= 32'hf50622a8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c8; din <= 32'h9b653efc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h158; din <= 32'hd1a77e40;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a4; din <= 32'h6872fa9c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d1; din <= 32'h105a513f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h340; din <= 32'h809540b4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15b; din <= 32'h6f7c39a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f6; din <= 32'hd08ff797;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cb; din <= 32'h8601f4d8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h398; din <= 32'he9ad99de;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13f; din <= 32'h3fe3412b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a7; din <= 32'h5c2369b7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e4; din <= 32'haf6037b0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32c; din <= 32'hac01dc64;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13e; din <= 32'heec8ac90;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d1; din <= 32'h8d611e76;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h056; din <= 32'hf3523bc8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3db; din <= 32'h1f49b003;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d3; din <= 32'h55865ea6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22e; din <= 32'h73f5a908;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03a; din <= 32'h0364e900;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a2; din <= 32'h5425e3ab;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h195; din <= 32'h80bf0957;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d3; din <= 32'h9e8eadfd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h071; din <= 32'haad36379;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a6; din <= 32'h089b5ad4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17b; din <= 32'hc824f1f5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e6; din <= 32'h120dd6e2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h001; din <= 32'h6f39db6b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a1; din <= 32'h64c13466;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ec; din <= 32'h62520c51;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26c; din <= 32'h7b443690;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03b; din <= 32'ha6f255e6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a7; din <= 32'hc38ee59a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h106; din <= 32'h056a6158;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h245; din <= 32'h71f1ee27;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h084; din <= 32'hdf01aadc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h329; din <= 32'hfa647f54;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h121; din <= 32'h603100a8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e7; din <= 32'hab50e506;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c4; din <= 32'hc97dae75;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c3; din <= 32'h1f029620;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1be; din <= 32'hea8075e4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a8; din <= 32'h2d32922a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00f; din <= 32'h3c421ed7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3df; din <= 32'hfd66101b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h127; din <= 32'hb20fd26b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cb; din <= 32'h15189422;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0af; din <= 32'h60ee0983;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37e; din <= 32'h5e4c8245;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16d; din <= 32'hbf8cd2e6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29e; din <= 32'hca829d83;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e9; din <= 32'hbaa4191e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38f; din <= 32'h253a3c68;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h126; din <= 32'hcbc51ddd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f0; din <= 32'h1d827e13;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h030; din <= 32'h94d646a5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f0; din <= 32'h1210113e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h133; din <= 32'h10f1ed92;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2be; din <= 32'h163cfa30;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0af; din <= 32'h02158334;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39a; din <= 32'h81b5935a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10b; din <= 32'h71aae53b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21c; din <= 32'h98ec667b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05d; din <= 32'h68131cf1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h305; din <= 32'haea1e763;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h128; din <= 32'h76c85ed5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2aa; din <= 32'h9bd3efd7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h010; din <= 32'h06174116;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f1; din <= 32'hc04950d9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c3; din <= 32'h67b445e8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d1; din <= 32'hc162667d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h077; din <= 32'hf547aa8c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h347; din <= 32'hc0d82713;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h125; din <= 32'he77914a1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h285; din <= 32'h5b13d96a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e4; din <= 32'hec2045c6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b4; din <= 32'h3c0da46a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h135; din <= 32'h1c7da340;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ec; din <= 32'hdcdff194;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a8; din <= 32'h2a8940b0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39b; din <= 32'h1e940dec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bf; din <= 32'h1dfb8da1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22d; din <= 32'h25cccb2e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08b; din <= 32'h12999787;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e9; din <= 32'h8a2d0283;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h180; din <= 32'hf7769eed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e8; din <= 32'hfc698eb2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d4; din <= 32'haa3f6f84;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h392; din <= 32'h869fce31;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13a; din <= 32'h30dfddc4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h269; din <= 32'hec427bb0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h003; din <= 32'h05c62e19;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32b; din <= 32'hfb0696b6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ce; din <= 32'hebef2ffb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23d; din <= 32'h56cb55b2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c4; din <= 32'hf3bc552a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d8; din <= 32'h854e3fb6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ae; din <= 32'hd68e62c7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d0; din <= 32'h04fd8a9c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h049; din <= 32'ha7a9e28c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ea; din <= 32'hde3b71a4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11e; din <= 32'h9473f81c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f0; din <= 32'h38a80650;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h014; din <= 32'hdc4b5a47;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h348; din <= 32'hfc6fda01;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f6; din <= 32'hcfdc349a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22a; din <= 32'h31e2ee60;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h062; din <= 32'ha07b6c05;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h363; din <= 32'h8bdc3601;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c9; din <= 32'h8d8e9a4e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ac; din <= 32'h4c2e0b0a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08e; din <= 32'h1c4ed579;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32c; din <= 32'h15098584;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10a; din <= 32'h49fdabf6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b5; din <= 32'h7bcee741;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d6; din <= 32'hc2f3f306;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33c; din <= 32'h267280dd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ce; din <= 32'hbd90b712;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h262; din <= 32'hf500b125;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c0; din <= 32'h07c6244a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h338; din <= 32'hde79cb25;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13f; din <= 32'h62651977;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ec; din <= 32'h7c6006d2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h098; din <= 32'h829d0829;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h314; din <= 32'hf09ee898;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10b; din <= 32'h45388ce2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20e; din <= 32'h1fcf7cc0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fc; din <= 32'h7d7e0575;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h369; din <= 32'h5f56dc69;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d2; din <= 32'h92992ff3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h291; din <= 32'h32c93e3a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a8; din <= 32'hd456678f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h329; din <= 32'hcc0d0f2c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18e; din <= 32'h72a7b320;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29b; din <= 32'h0455c0c6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h008; din <= 32'h880db2d1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h393; din <= 32'h4c73295e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e9; din <= 32'h6d9051da;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h259; din <= 32'hab86013d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02e; din <= 32'he035cd29;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h342; din <= 32'h149e63a7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13c; din <= 32'h3b89bbb7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2fe; din <= 32'h0608c929;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09d; din <= 32'h04edee8b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h316; din <= 32'h5e8a51b4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ab; din <= 32'hdf1024b0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e3; din <= 32'h27f494ef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h088; din <= 32'hcc18f91e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33a; din <= 32'hed9ea1e9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16c; din <= 32'h4dad0d2b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h250; din <= 32'h58783c03;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d1; din <= 32'h8b52443d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h365; din <= 32'h229999ad;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a2; din <= 32'hf2fc365c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26b; din <= 32'he0fbbf12;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fc; din <= 32'h64bc1475;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f3; din <= 32'h2ccf3d42;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c9; din <= 32'hc735d632;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27d; din <= 32'h13745351;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03b; din <= 32'h2abf03d2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h338; din <= 32'he1bbfca3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17f; din <= 32'h03d91034;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a7; din <= 32'hc9f2cce7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h070; din <= 32'h9f3a0dbc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d8; din <= 32'h1ffed833;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h188; din <= 32'hcb360808;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h291; din <= 32'hfe801c4a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h070; din <= 32'h2ca2bbc9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38c; din <= 32'he77bc5e3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h148; din <= 32'h5fe7453a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26c; din <= 32'h80dcb333;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e2; din <= 32'ha5c5c464;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c7; din <= 32'h386aa4a2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13e; din <= 32'heb058e45;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h283; din <= 32'h1821ac02;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a1; din <= 32'h585fad3b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32c; din <= 32'h6234f9e8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h108; din <= 32'h21e761eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h288; din <= 32'hcf58c36c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fd; din <= 32'h104ab3d6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f7; din <= 32'h5a881424;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13e; din <= 32'h6e83a783;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ab; din <= 32'h3605fde3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d8; din <= 32'h7d3e4d5c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cb; din <= 32'h4c4e7e34;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h167; din <= 32'h821c2bc5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a7; din <= 32'h3bc9fbe2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0dc; din <= 32'he77fb785;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ef; din <= 32'hb359a454;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12f; din <= 32'h99be1a3e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h251; din <= 32'hd87713e5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h088; din <= 32'h8004a634;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d3; din <= 32'h77354dee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18a; din <= 32'h821d64ce;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h281; din <= 32'hba61b206;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fe; din <= 32'h6d8aa9ab;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32e; din <= 32'hfdfc2fbf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h192; din <= 32'h8492e939;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d0; din <= 32'hd5e65816;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a8; din <= 32'h557a8b28;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36c; din <= 32'h07c86d1e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e5; din <= 32'h9b01e6ed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h217; din <= 32'h85bdf8ca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c5; din <= 32'hd65c2a58;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ce; din <= 32'hbace02c2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h165; din <= 32'hc903ba73;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27e; din <= 32'h29354a83;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h053; din <= 32'ha932976f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31d; din <= 32'hbb3a23b6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cf; din <= 32'h72dfb536;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27a; din <= 32'he6bd2355;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a7; din <= 32'h004a3013;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f6; din <= 32'h45a246f7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1db; din <= 32'h1c329b65;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21b; din <= 32'h7df47e85;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03f; din <= 32'hc5ef538d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32f; din <= 32'h1a09966f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h169; din <= 32'h6af6e8a3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d7; din <= 32'h6ed5a774;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05f; din <= 32'h7eee573e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c7; din <= 32'h9a6bba8a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h184; din <= 32'h85d3d872;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27d; din <= 32'h1f9b23d5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e2; din <= 32'he295c038;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c8; din <= 32'h76dfd0d3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16c; din <= 32'h9246fca9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20f; din <= 32'h7ee4cea0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00a; din <= 32'he5c2bdf3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33d; din <= 32'h92994fde;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d4; din <= 32'h684fcf0e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h214; din <= 32'h5a3ff27f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f8; din <= 32'h2e8daa75;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h391; din <= 32'hc6f4f0c0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h166; din <= 32'h1d297576;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h281; din <= 32'hdbd66ee0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e4; din <= 32'h20c1efe0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d0; din <= 32'h6cc8738a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11d; din <= 32'h676296f3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2dd; din <= 32'h2daa130c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h050; din <= 32'hce7be123;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ee; din <= 32'h96dee588;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c2; din <= 32'h7b945756;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h252; din <= 32'h040beb3e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06e; din <= 32'h90d0dd42;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e4; din <= 32'h11bd3eb4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bf; din <= 32'h27213cab;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h274; din <= 32'hb2581cfd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h007; din <= 32'h6792aa08;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h397; din <= 32'h69f75573;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h126; din <= 32'h7b9d5243;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h285; din <= 32'hf0a2851e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h019; din <= 32'he219ce5a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h332; din <= 32'h37e5e5cc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h172; din <= 32'hf52316e6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h203; din <= 32'h678f9b21;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h013; din <= 32'hc327c5c0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fb; din <= 32'h581d48d8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1de; din <= 32'h6bc29651;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h293; din <= 32'h20b3a396;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h058; din <= 32'he742374c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c8; din <= 32'h298278fb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d7; din <= 32'h806fdb8d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h248; din <= 32'hdda7c99d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f2; din <= 32'h9322d46f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33c; din <= 32'h2936a3ad;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e8; din <= 32'h7f7a9346;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h285; din <= 32'h64c7eefe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h097; din <= 32'h92419d6f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h394; din <= 32'hc750fadf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10e; din <= 32'hf11faacb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24f; din <= 32'h6bc34865;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h098; din <= 32'h7d4bae8c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h390; din <= 32'h40503ee0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h115; din <= 32'h23b5a488;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2af; din <= 32'hb7737f2c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h083; din <= 32'hef951a0e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h361; din <= 32'h6dc94463;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13d; din <= 32'h35b4052d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b0; din <= 32'h1057c77b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h045; din <= 32'h5179ac44;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h336; din <= 32'h130662ac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h196; din <= 32'hfb9047b7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ad; din <= 32'h6f92c1fe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h096; din <= 32'h242b258d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e6; din <= 32'hcef83dde;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h127; din <= 32'h3016934e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2aa; din <= 32'h87d916c1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e0; din <= 32'h918b6b16;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f2; din <= 32'h48fa599d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h109; din <= 32'hc77e4d93;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23c; din <= 32'h61d8352f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h078; din <= 32'h9709df62;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fe; din <= 32'h893c7cb8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fd; din <= 32'h3eabed6d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h260; din <= 32'h041c8d9a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04e; din <= 32'h3a678b9d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h355; din <= 32'h65f84cf1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1df; din <= 32'hebf49a72;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h261; din <= 32'hb2f4a827;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0be; din <= 32'h929da2d8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h308; din <= 32'h86c578af;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ed; din <= 32'h3ae4d1da;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28b; din <= 32'h71d5f103;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c2; din <= 32'h483b3ec4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h373; din <= 32'hdcd20046;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10e; din <= 32'hcdd4bb9d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h239; din <= 32'h7ead3b6d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07b; din <= 32'hc36fee67;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h355; din <= 32'h9b98be96;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f2; din <= 32'h228f31f7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23d; din <= 32'h235b38c8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e8; din <= 32'h966bd9f9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h343; din <= 32'hba31c376;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b9; din <= 32'h80eb896d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h234; din <= 32'h14606825;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04f; din <= 32'h8820b02d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37f; din <= 32'h54a89f46;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fa; din <= 32'h414e331f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h228; din <= 32'he5b86229;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h073; din <= 32'hfa5d3e8c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35a; din <= 32'h14b43a2a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ab; din <= 32'hb5a43767;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21b; din <= 32'hb708397f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h077; din <= 32'h3c15cec3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34b; din <= 32'hea58687e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h197; din <= 32'h78a61992;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h277; din <= 32'h6112f2e4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ba; din <= 32'hdc1b2a06;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30e; din <= 32'h5f725313;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h165; din <= 32'hdb4fea5a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22a; din <= 32'h4fd5b3f3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d1; din <= 32'h0337dc44;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39e; din <= 32'hfd722c5f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14c; din <= 32'had744cd3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21b; din <= 32'h27c19e84;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c6; din <= 32'h63130428;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fe; din <= 32'h71498d58;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h173; din <= 32'hf3b144e7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c3; din <= 32'hc7fee970;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c5; din <= 32'hbc3e4eb0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h372; din <= 32'h78055fa7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d3; din <= 32'hd851d37b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h219; din <= 32'h9f3813e0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b6; din <= 32'hb2cd849c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h366; din <= 32'hf610181e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b2; din <= 32'hbb3acf65;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h267; din <= 32'h76a3d754;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01e; din <= 32'h8adb0722;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h324; din <= 32'h6fed3965;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h110; din <= 32'h9be49032;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27e; din <= 32'hbb5a8dce;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01f; din <= 32'hf23c8808;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h394; din <= 32'h0a583a35;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h163; din <= 32'hbc6f3374;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h240; din <= 32'h07403a5a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c6; din <= 32'h1155fef4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h332; din <= 32'h45dd933f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h175; din <= 32'h56679a79;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h213; din <= 32'h39397d64;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h032; din <= 32'hb5725391;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h390; din <= 32'hcf4bb5c0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h116; din <= 32'h9aefa186;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h283; din <= 32'h31382496;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a5; din <= 32'h32f777eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d5; din <= 32'hf04cbec4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18f; din <= 32'hd98f7d04;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e9; din <= 32'he5e50b0e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h077; din <= 32'h6aa59fe1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bd; din <= 32'h89adc337;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16f; din <= 32'h5a84a3f8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h271; din <= 32'h69f5000e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09a; din <= 32'hfef6a625;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f5; din <= 32'hba038b56;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d0; din <= 32'h39bb253b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22a; din <= 32'hd6636300;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e1; din <= 32'h77510435;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3dd; din <= 32'h73fda743;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ad; din <= 32'h72e028e5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h228; din <= 32'h53565d30;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d8; din <= 32'h551ed5d5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h395; din <= 32'hcb28418c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h158; din <= 32'h29ee99c6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h249; din <= 32'h03f84c07;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01b; din <= 32'h0336c518;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h397; din <= 32'h6145cc78;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h122; din <= 32'h59f06ef1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21c; din <= 32'hec06c91a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h044; din <= 32'hdfe4cbd7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37a; din <= 32'hd1403cd9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10c; din <= 32'h9c07e092;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h227; din <= 32'hc62a7990;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05b; din <= 32'hcddf02e8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f8; din <= 32'h266401d6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h105; din <= 32'h2502fc4b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h212; din <= 32'h3422e0a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h088; din <= 32'h2b7793db;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c8; din <= 32'h5b637e6e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f7; din <= 32'h8fd7e9e2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h290; din <= 32'h24c65b4b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07a; din <= 32'h1fec9c4b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h314; din <= 32'h155e8bc3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h183; din <= 32'h85c1cc26;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29a; din <= 32'he7d2c764;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00c; din <= 32'hcdf18bd2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h396; din <= 32'h85f7eb7a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ab; din <= 32'hfcb0c40b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h284; din <= 32'h73fbfba5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0de; din <= 32'he4f8f3ac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cc; din <= 32'h3eabb7ae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1df; din <= 32'h6ab64441;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28e; din <= 32'hc940d751;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h079; din <= 32'h48b73875;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34a; din <= 32'hbee43262;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18d; din <= 32'hde89c21a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h275; din <= 32'hf155d8c1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h062; din <= 32'h4aab1994;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h319; din <= 32'he50b35e2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cc; din <= 32'h5d887ab3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ea; din <= 32'hfe0023c7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h072; din <= 32'hbd08b43e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h382; din <= 32'h1ce12967;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17c; din <= 32'h39bf769f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h219; din <= 32'hd2a89456;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h066; din <= 32'hac6f9188;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ca; din <= 32'h4a153357;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b3; din <= 32'h22437070;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h279; din <= 32'h074f600e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h058; din <= 32'h519e495f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h388; din <= 32'hae5405a8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16a; din <= 32'h0f3b374f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e3; din <= 32'h212f66c0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e6; din <= 32'hdd75cfb8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30c; din <= 32'h6df71144;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15e; din <= 32'hb4a60e0a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23d; din <= 32'hc49e9247;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08f; din <= 32'h4c308c14;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a4; din <= 32'he4fdfdcc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h165; din <= 32'h54e922fd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h266; din <= 32'hf6b5b41e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05b; din <= 32'hc1b627e0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f8; din <= 32'haa3f58f9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h117; din <= 32'h235917a3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27e; din <= 32'hbb405824;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0eb; din <= 32'h95ed9643;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h314; din <= 32'hf4d9b75a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f8; din <= 32'h2c2d10aa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ab; din <= 32'h99668a18;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h043; din <= 32'hfc0beea0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d7; din <= 32'h14e65919;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h136; din <= 32'h7fa5a5dc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f8; din <= 32'ha3386ea7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a7; din <= 32'h33bd8aae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h357; din <= 32'had9e0569;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h129; din <= 32'hc30fd932;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a1; din <= 32'hd0c526c6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h028; din <= 32'hb9ad217f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e3; din <= 32'ha71a196e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f6; din <= 32'h37fe6397;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e4; din <= 32'hc5af50d4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h013; din <= 32'hed01b777;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c4; din <= 32'h9284923f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ad; din <= 32'h3bcd5cf2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h277; din <= 32'h7c3bb743;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h006; din <= 32'h76a38c5d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a9; din <= 32'hf7ec9708;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h178; din <= 32'hd3ba2dac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e4; din <= 32'h9ec6298b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02c; din <= 32'hb85aca79;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ed; din <= 32'h7d95e484;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f9; din <= 32'h95cce965;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bb; din <= 32'hf9c4895b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c7; din <= 32'hfe084cec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b3; din <= 32'h082a6d4e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cb; din <= 32'h56f0c952;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f2; din <= 32'h1a65c7b1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06c; din <= 32'h64c1d9c5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b7; din <= 32'h089db854;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d7; din <= 32'hc92420b7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a6; din <= 32'hc7f7efaa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02b; din <= 32'h103035cf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32d; din <= 32'he32bf11c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fc; din <= 32'h5cf677af;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28c; din <= 32'ha5fb55bf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h078; din <= 32'h86ac803b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h393; din <= 32'h5aef34d2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14b; din <= 32'he9c8f333;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20d; din <= 32'h1111f860;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06a; din <= 32'h25c81829;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h334; din <= 32'h6cd96293;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h194; din <= 32'hcb810100;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27d; din <= 32'hcb13b9df;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01d; din <= 32'h7037d31a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h395; din <= 32'h498c3d7d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h177; din <= 32'hd7c8bc55;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h210; din <= 32'h2e3cd420;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08c; din <= 32'h0e16011f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h385; din <= 32'h260af13e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d9; din <= 32'haf36efe9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h277; din <= 32'h297d783f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h033; din <= 32'h09c1341d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cd; din <= 32'heb938b52;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h141; din <= 32'h861bcd1c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h209; din <= 32'hf8db64da;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c0; din <= 32'h34fc3a87;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h377; din <= 32'h3d85748b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1df; din <= 32'hb459b9fc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h263; din <= 32'h3ce6b4ba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07b; din <= 32'h0ece5adb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h344; din <= 32'h5ec5e57d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ba; din <= 32'h5767db54;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h298; din <= 32'h3c68e4cc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07c; din <= 32'h11df6247;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h352; din <= 32'h8209d65e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cc; din <= 32'h2eeaabce;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2eb; din <= 32'h5aec71a7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h082; din <= 32'h51a2d4a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32e; din <= 32'h83be072b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h111; din <= 32'h1b73f289;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h239; din <= 32'h35cd9f6b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ad; din <= 32'he2ff05c9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h317; din <= 32'h29a0e486;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1eb; din <= 32'hec8c335c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cf; din <= 32'h0f1b640e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c7; din <= 32'h60a0492e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a9; din <= 32'h04e73878;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h122; din <= 32'ha0b2a7c6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c9; din <= 32'h84f9dd1a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e8; din <= 32'hf1bdcda0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a6; din <= 32'h3aa82292;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b1; din <= 32'h89eeda77;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bf; din <= 32'h3bc61afd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c3; din <= 32'h04048a85;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d1; din <= 32'h274d4832;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h112; din <= 32'h19c93111;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d1; din <= 32'h2b6167a1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cc; din <= 32'hf10a05f4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37f; din <= 32'hdc9ede6c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bf; din <= 32'ha38c20b0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h209; din <= 32'h38f1d03d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h060; din <= 32'h52671507;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38a; din <= 32'he3251430;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10a; din <= 32'hac3d8f0c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2eb; din <= 32'h45acaff8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h033; din <= 32'h32f62d68;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h320; din <= 32'h608ee225;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ac; din <= 32'h208e458a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h273; din <= 32'hd41b5cf2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02d; din <= 32'h8d04fea1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33d; din <= 32'h06a370e3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12b; din <= 32'he7607b84;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h289; din <= 32'hf7f3ab81;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f2; din <= 32'hbe18f5be;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h396; din <= 32'h28c6df0e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h160; din <= 32'h6422ce96;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24c; din <= 32'h5b32d0ca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05e; din <= 32'h7876bec8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h327; din <= 32'h6e36930b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h182; din <= 32'h0bf36199;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h214; din <= 32'h52ccf0bd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h084; din <= 32'h676486fd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cc; din <= 32'h52aadd19;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h111; din <= 32'h0d9ceea1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24f; din <= 32'hc63c330f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d4; din <= 32'h712ac8d2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c6; din <= 32'he5d292d6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h118; din <= 32'hf144da97;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e6; din <= 32'h41d4e271;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h082; din <= 32'hb610ec0e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h332; din <= 32'ha07a0efc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h190; din <= 32'h0de9ff36;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h270; din <= 32'h25bd7782;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h027; din <= 32'he2b7b27a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a0; din <= 32'h9ec0bde8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h123; din <= 32'h95fb9123;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27b; din <= 32'h0f5abe76;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h022; din <= 32'h4ec41279;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b1; din <= 32'h1051faa7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18d; din <= 32'h4d17a8ee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29d; din <= 32'h6be24aea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h098; din <= 32'h9416df51;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34f; din <= 32'h5d5fadef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h167; din <= 32'heb913d16;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a8; din <= 32'hd98c67b5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h082; din <= 32'hb1e685b0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34b; din <= 32'h4eafcd98;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h165; din <= 32'h34a40f7c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e8; din <= 32'h97b47d6a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09e; din <= 32'h73b18036;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h386; din <= 32'h91c20eee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bb; din <= 32'h3bc57d2d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h276; din <= 32'h8d6620e5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h008; din <= 32'h9e92a667;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33a; din <= 32'h340bac94;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ba; din <= 32'h9c8fcb33;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e2; din <= 32'h0b1db824;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h064; din <= 32'h7bcf97e1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38a; din <= 32'hafcbcbd8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d7; din <= 32'h52f0168f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h287; din <= 32'h196a4707;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05e; din <= 32'h80a37a34;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f9; din <= 32'h9bab9a7e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h174; din <= 32'h890d58ea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h206; din <= 32'hfbe6a9ff;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f6; din <= 32'h46b5e33b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h325; din <= 32'hd85ba608;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a8; din <= 32'h714d7280;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h201; din <= 32'h45437062;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h089; din <= 32'hf88a85d2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39b; din <= 32'h85136b4b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a7; din <= 32'he5b1de29;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22e; din <= 32'h04ff9889;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h037; din <= 32'h9abc9e79;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3eb; din <= 32'h66959e81;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cf; din <= 32'he82c5ff3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h233; din <= 32'h93b79828;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b5; din <= 32'hd3e780ef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3dc; din <= 32'h817c6fda;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14b; din <= 32'hcc567c42;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h240; din <= 32'h8ca2cffb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ca; din <= 32'h4f98b627;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30f; din <= 32'hee3b6b36;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19b; din <= 32'hfaf31e0c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h254; din <= 32'h57abf690;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d2; din <= 32'h4d8f7ee1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h391; din <= 32'h92bd61e7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h175; din <= 32'h45a9449b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e2; din <= 32'h46e06ed2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f6; din <= 32'h39c3ea9d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h387; din <= 32'h608444c4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10f; din <= 32'hdcfb9d28;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cc; din <= 32'hd7b2557a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ae; din <= 32'hc1b8c86d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h348; din <= 32'hf742dbd4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15b; din <= 32'h09d22a9d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22f; din <= 32'h87987209;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e3; din <= 32'h34cf1fff;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a8; din <= 32'h8df71700;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h149; din <= 32'h47958aad;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h237; din <= 32'h278a6bda;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h003; din <= 32'h45a6b922;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h374; din <= 32'hdccdc260;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fe; din <= 32'hf9eda88b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ec; din <= 32'hc9fc8aee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c9; din <= 32'haa3f77cb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h340; din <= 32'h8de5ae71;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f6; din <= 32'hbb4e063f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24e; din <= 32'h9deaefe5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h010; din <= 32'h97cb484b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a3; din <= 32'hc08ce807;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e7; din <= 32'hb336b63f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h270; din <= 32'hf1bc36dd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05b; din <= 32'h8cf7111a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h353; din <= 32'h7c35c774;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cb; din <= 32'h9c0cd630;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h270; din <= 32'hc448f832;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h069; din <= 32'h746fa068;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h363; din <= 32'h4284b9ce;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16e; din <= 32'hc1340a04;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c8; din <= 32'h74e406ac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bc; din <= 32'hfef523d0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fb; din <= 32'hf4314c5e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d5; din <= 32'he88d66a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25f; din <= 32'h7eec57bd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h025; din <= 32'hee931a6d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cf; din <= 32'hfad1ec0e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15a; din <= 32'hc55aea50;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b4; din <= 32'h2211e9c1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h077; din <= 32'h6fe049f5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ea; din <= 32'ha8c5345f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h137; din <= 32'h7171fc7f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25e; din <= 32'h4d399089;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09c; din <= 32'hcd9e0f92;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h315; din <= 32'hb699cff1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f6; din <= 32'h76a9ea9a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h255; din <= 32'h3d3c0a7a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h043; din <= 32'hb867f347;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3aa; din <= 32'ha6a4321f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bf; din <= 32'h1b1d43ca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h264; din <= 32'h9ba43e54;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h082; din <= 32'h72d45776;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h351; din <= 32'hf35cbad7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15a; din <= 32'h65aafb7e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f3; din <= 32'hed15ff05;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08b; din <= 32'he5ff2c5e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h365; din <= 32'hc5ac6c1b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h121; din <= 32'h0a7574e1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h286; din <= 32'h3025bac8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fa; din <= 32'h1e501b77;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h377; din <= 32'h520c20e0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h185; din <= 32'hb4f49eae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a6; din <= 32'hc422e393;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c6; din <= 32'h073e4e08;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38e; din <= 32'h809718ec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c4; din <= 32'hf80ba61f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22f; din <= 32'h8076ad31;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bf; din <= 32'h09ce01a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h367; din <= 32'h1d4f5bb7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h149; din <= 32'h8fa84a77;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27f; din <= 32'h19fe7ab5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h082; din <= 32'ha980493c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d8; din <= 32'h1a129aab;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11b; din <= 32'h8cd08e8c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28c; din <= 32'h926e650b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04d; din <= 32'hf88c0aaf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39d; din <= 32'hec788878;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h119; din <= 32'hc751915e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e9; din <= 32'hed913241;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08b; din <= 32'h8fb9d3e0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h328; din <= 32'h48013c09;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d0; din <= 32'h1bba4a91;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21c; din <= 32'hc730bf6d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d1; din <= 32'h27251ae9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c6; din <= 32'h3d3f375c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h114; din <= 32'he7ba5459;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h284; din <= 32'ha8af85d5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h007; din <= 32'h1c2df1aa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h340; din <= 32'h7396eb9f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1da; din <= 32'haaeaa883;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a7; din <= 32'h48cd0374;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09a; din <= 32'h4bc57705;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32f; din <= 32'he27e3617;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d4; din <= 32'h1fbae6c9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27a; din <= 32'h55da7137;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h039; din <= 32'hfb0828d0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37f; din <= 32'h2b008826;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b0; din <= 32'h53ac8694;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2eb; din <= 32'h86f9fb0c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05e; din <= 32'h76ef6d15;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h313; din <= 32'ha4941a42;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a2; din <= 32'h194e3cc1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h228; din <= 32'h83542f43;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h014; din <= 32'hcaacffc6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d7; din <= 32'h79c6d99e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fd; din <= 32'ha0ba3a57;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23b; din <= 32'hef22f211;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a2; din <= 32'h28c86af7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ab; din <= 32'h2582324f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h140; din <= 32'h835218a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h276; din <= 32'he32f03e2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a1; din <= 32'hcb194db5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h326; din <= 32'h52c76d85;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10d; din <= 32'h2e9f3c78;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22d; din <= 32'hf4914a08;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0af; din <= 32'hc2b13373;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h318; din <= 32'h082a2f29;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d8; din <= 32'hfaf2367b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c3; din <= 32'h0e344131;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f6; din <= 32'h1216ac39;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30f; din <= 32'h08a83ebe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c7; din <= 32'h2c6e54d6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e1; din <= 32'h2da4eae8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fe; din <= 32'h0132b0b4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h342; din <= 32'hdf8e976d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e5; din <= 32'h74cf3805;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a9; din <= 32'h9487ad7a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bb; din <= 32'ha40b0257;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ea; din <= 32'hf7c8c198;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18c; din <= 32'h787188f8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24e; din <= 32'h50aa4b38;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c5; din <= 32'h28a3b600;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a8; din <= 32'hb2646699;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h185; din <= 32'h99342c54;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26e; din <= 32'hbcfe2d96;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02e; din <= 32'hb42613c3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37f; din <= 32'h40f145ac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13b; din <= 32'ha1e5bbca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h246; din <= 32'hb34ba26e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04e; din <= 32'hc8b5ed5a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b6; din <= 32'h7d000be6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1db; din <= 32'h0fccd7da;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h298; din <= 32'hcda7a356;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h004; din <= 32'h83b129cd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a3; din <= 32'h653ca2cd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h120; din <= 32'h6ff71f0e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23f; din <= 32'h80a60962;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h063; din <= 32'heceb9a4c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fc; din <= 32'he1d680eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17e; din <= 32'h93cdb56a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f7; din <= 32'h122daaa5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h009; din <= 32'h457b43f1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e7; din <= 32'h05bbf21b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h177; din <= 32'h49c9f06e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d3; din <= 32'h4ab71c66;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03b; din <= 32'h862c5655;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39d; din <= 32'h27047bdd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cc; din <= 32'h075495ba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b1; din <= 32'h33c2fbf4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07b; din <= 32'ha1488f83;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fe; din <= 32'h92661b7d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bd; din <= 32'hf1c936cf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27e; din <= 32'h59926876;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ec; din <= 32'hec469526;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h307; din <= 32'hf886f267;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e0; din <= 32'h056bfbe6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2de; din <= 32'hf6499cf3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h019; din <= 32'h5724a618;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33f; din <= 32'h1f1dc796;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16d; din <= 32'h435b129a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23e; din <= 32'h5666ac3f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h058; din <= 32'hd57bf316;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h312; din <= 32'hdacc3b52;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h147; din <= 32'hddc168d9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29f; din <= 32'hb811d528;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a7; din <= 32'hffd40925;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h309; din <= 32'hcae8d54a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h140; din <= 32'h3ee53c6d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26d; din <= 32'h902d4d58;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03c; din <= 32'hbb121509;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32d; din <= 32'h2c7af735;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12b; din <= 32'h23750d90;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e5; din <= 32'h6a37e53c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h057; din <= 32'hda59dd29;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32b; din <= 32'hc66a1e97;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ee; din <= 32'h177e3ecf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c4; din <= 32'hb4df7ed8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h059; din <= 32'h4bfd1559;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d3; din <= 32'hf674ad8e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16d; din <= 32'h4fb4f75c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h210; din <= 32'h419d00ea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0aa; din <= 32'h079020fc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h329; din <= 32'hc18bac53;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ea; din <= 32'h164e9298;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h297; din <= 32'hc538ea87;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a6; din <= 32'h79fb8fdd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h363; din <= 32'h5b266047;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h100; din <= 32'h5ab5cc70;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h215; din <= 32'hfb74e860;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cd; din <= 32'h031562d6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h356; din <= 32'h246eb2fa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h194; din <= 32'h7d8b7548;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h234; din <= 32'h5c19ac9a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h019; din <= 32'h16463616;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h301; din <= 32'h9d3b0072;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h198; din <= 32'ha8b24e2d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24b; din <= 32'hc6aa6aca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a3; din <= 32'h78a00ca4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h390; din <= 32'h441e359c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d7; din <= 32'h6dceb9e8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h223; din <= 32'hf031eb80;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h001; din <= 32'h42d4cc55;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ef; din <= 32'h7887762f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18b; din <= 32'hb6254f23;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b4; din <= 32'h4966c501;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h079; din <= 32'h0b580aa7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e7; din <= 32'hd7b09da9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h154; din <= 32'h3ea5b091;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ba; din <= 32'h53ba17e3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h072; din <= 32'h7f9f2556;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c1; din <= 32'h69e757a2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16f; din <= 32'h7d576f5d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h220; din <= 32'h7b428c66;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d1; din <= 32'h6b819056;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h395; din <= 32'h02aeade8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e7; din <= 32'h5cf09272;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28d; din <= 32'hb616abea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f3; din <= 32'h28c28220;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30a; din <= 32'h3be199d0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h126; din <= 32'hfc3ad404;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b0; din <= 32'h9f5caa17;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04f; din <= 32'hbd9e6a9c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32d; din <= 32'h847271d3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17b; din <= 32'hbe85e2c6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a8; din <= 32'hf00be967;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ee; din <= 32'hcbcddae4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h352; din <= 32'h732bb6ab;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h157; din <= 32'h9ee2fb0d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b9; din <= 32'h7eb00c7b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h085; din <= 32'h69b1c57b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3df; din <= 32'hf5fbcec2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h111; din <= 32'h893e2bbf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2de; din <= 32'he3a9005d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h049; din <= 32'h0afaa2ac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h387; din <= 32'hfccb7ba0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a8; din <= 32'ha0b6a413;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c3; din <= 32'h6b825d47;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h003; din <= 32'h368642d7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bb; din <= 32'h78d0b892;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14f; din <= 32'h04cee693;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h205; din <= 32'hf0fe86b5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h058; din <= 32'h532b9289;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h382; din <= 32'h3771213b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12b; din <= 32'hfe2bb1f7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bb; din <= 32'heb0b6c50;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b1; din <= 32'h642e3b4a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h307; din <= 32'h33698c37;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16c; din <= 32'h024db6de;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h271; din <= 32'h98ae9c80;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h078; din <= 32'ha4e9e6ae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fc; din <= 32'hcabb4d19;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a9; din <= 32'h00f693fa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26f; din <= 32'h03791279;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06e; din <= 32'hb82d212e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35a; din <= 32'hea75ea17;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h146; din <= 32'h07fdbe2e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h223; din <= 32'h6a78a6be;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b2; din <= 32'he661655c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34a; din <= 32'h907f6d0b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c1; din <= 32'hd354b2d5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29d; din <= 32'ha3cbc494;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d6; din <= 32'hc6a73204;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h323; din <= 32'hde67dc39;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h103; din <= 32'h1859b805;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h211; din <= 32'ha8a7e3d5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h096; din <= 32'hd924013e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38d; din <= 32'h728a91cd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17e; din <= 32'h0cf7f337;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h257; din <= 32'h8ee4b91d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fa; din <= 32'h0d31a88d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h305; din <= 32'hc1aac481;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h135; din <= 32'hb560d92a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20a; din <= 32'ha6165e5a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h094; din <= 32'h7ffbd8f7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h321; din <= 32'h1b9e4c5d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h113; din <= 32'h4649bcf0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f5; din <= 32'h96777382;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h056; din <= 32'h4c684903;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34a; din <= 32'h4fc94a09;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c0; din <= 32'h60e4f986;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h274; din <= 32'hecd80ffd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h028; din <= 32'h306e3577;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30c; din <= 32'h14fd17cb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h164; din <= 32'h89770b41;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cc; din <= 32'h49fae24c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e4; din <= 32'hcd283643;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f0; din <= 32'hfaabb64a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14e; din <= 32'h780777ee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h202; din <= 32'h81d25c2e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a7; din <= 32'h5905ee98;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39a; din <= 32'h44c637b2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h175; din <= 32'h06880bf3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h242; din <= 32'h568a22b3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03f; din <= 32'hefcb71fd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d6; din <= 32'h5b49fcb8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h179; din <= 32'h559ea3ea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25b; din <= 32'h7114e5dd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05c; din <= 32'hb4386164;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3db; din <= 32'hb16aaabe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c0; din <= 32'h599b7094;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cb; din <= 32'hf4c8fde2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ab; din <= 32'hd64d0968;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ef; din <= 32'hf553e0a1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d5; din <= 32'hc3eaa0d2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h224; din <= 32'h39b0630a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cc; din <= 32'h96b08134;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h334; din <= 32'h8b0268df;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c0; din <= 32'h24baf923;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25f; din <= 32'hd10a67dc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01e; din <= 32'h55bc9519;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38f; din <= 32'hd20911e1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h195; din <= 32'h038dd32d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20a; din <= 32'h530ad4b8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ae; din <= 32'h1f37ad26;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h392; din <= 32'hbda1ca20;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c3; din <= 32'h6f31c6d8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26e; din <= 32'h281ec149;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h066; din <= 32'h2260c633;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34d; din <= 32'h60e1bce8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ac; din <= 32'h98001268;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b4; din <= 32'h2028d5a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bb; din <= 32'h514a30b9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h313; din <= 32'hfa9684ab;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17f; din <= 32'hc58df5aa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h253; din <= 32'h11cd5300;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h024; din <= 32'hb5ac6344;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h377; din <= 32'hb253e343;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h110; din <= 32'h4439ed93;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21b; din <= 32'h4a1cac26;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h016; din <= 32'h934ca534;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h355; din <= 32'he050c200;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16a; din <= 32'h326da00e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h273; din <= 32'h4bd373d3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cd; din <= 32'hb5e1b861;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31a; din <= 32'h1600c62e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ab; din <= 32'h0daf8fbd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20f; din <= 32'h4c55ac95;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h060; din <= 32'h91d53798;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34d; din <= 32'h28d46b7e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h174; din <= 32'he604aa41;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25d; din <= 32'h3450b928;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h040; din <= 32'h0d631e9e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f3; din <= 32'ha6852fcf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h115; din <= 32'ha85613f8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ed; din <= 32'h5fed3032;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f5; din <= 32'h742d7e27;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e2; din <= 32'h08a9463b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h130; din <= 32'hb3723371;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21b; din <= 32'h408d9f37;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ec; din <= 32'h5a1ad941;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h343; din <= 32'h7a05ec04;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e4; din <= 32'h86b53705;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h295; din <= 32'h8d25fbea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h072; din <= 32'h30c4a0dd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b1; din <= 32'he1533d8e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13c; din <= 32'h4dd3c6f8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h254; din <= 32'h9280c827;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fa; din <= 32'h0b7504f6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b4; din <= 32'h8c2c18f8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h123; din <= 32'h3a65366c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2df; din <= 32'h5f23a6af;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c8; din <= 32'h25398ef5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d6; din <= 32'h24279760;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19e; din <= 32'h037d62c0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c5; din <= 32'h800f3036;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00f; din <= 32'hd6acb9eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39a; din <= 32'h0c33080f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16b; din <= 32'hb1a87e1b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h256; din <= 32'hef949cde;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h010; din <= 32'h84a538ae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h360; din <= 32'hfc240d72;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h185; din <= 32'he29e6ed4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21c; din <= 32'h6c1d80eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03f; din <= 32'h79c8326d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31a; din <= 32'hf1225e95;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11d; din <= 32'h2bf64255;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2db; din <= 32'h0629f585;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h093; din <= 32'h4373f1ab;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3de; din <= 32'h61083974;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19b; din <= 32'h433314b0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2eb; din <= 32'h45934ef1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c1; din <= 32'h5dfc59de;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bb; din <= 32'h5f62e799;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h186; din <= 32'h5f647fa3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h250; din <= 32'h53d6b10e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h052; din <= 32'hd782c57e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d3; din <= 32'h1c12c841;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f1; din <= 32'hf8556f5f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ee; din <= 32'he3413c8a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h079; din <= 32'h23abaa9a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h306; din <= 32'h418847eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h114; din <= 32'hf6323951;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bd; din <= 32'hd4d68830;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h069; din <= 32'h78ccf50c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38f; din <= 32'h0b2d5208;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16c; din <= 32'h384f9da2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ec; din <= 32'hca025b0c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h049; din <= 32'h0f8ef202;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ec; din <= 32'hdbed1d5f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d6; din <= 32'hc1d5d61e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25c; din <= 32'h631a6f17;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f2; din <= 32'h80a69fb3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h342; din <= 32'h140a91b8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13d; din <= 32'hf3d5ee42;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d1; din <= 32'hfbb67d38;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b6; din <= 32'he7af15c6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h310; din <= 32'hb3fb3e1e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d1; din <= 32'h3c76dc08;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h210; din <= 32'h501b66b4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d7; din <= 32'h109c89e2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37f; din <= 32'h2275085a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13e; din <= 32'h5e3e6c68;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b4; din <= 32'hc44255f5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h040; din <= 32'h5516e8da;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h380; din <= 32'h665c16d1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h166; din <= 32'hb4522a47;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h235; din <= 32'h2af89c10;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c8; din <= 32'ha248bae7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b5; din <= 32'hc815aa35;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h122; din <= 32'h2588ae3b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d5; din <= 32'he721a1f5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e4; din <= 32'hca889340;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35d; din <= 32'ha2cfcfcb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d9; din <= 32'h0c0bc2e8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d0; din <= 32'h56f7ab85;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b4; din <= 32'hd3c00c7a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h337; din <= 32'hf070a3b7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h176; din <= 32'hfde05b92;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h231; din <= 32'hbb6745ce;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e4; din <= 32'h60a64a9c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35f; din <= 32'h6ad3c68e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cb; din <= 32'hbfab7d32;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27e; din <= 32'hd1767636;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f7; din <= 32'h7ec8e7c6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ab; din <= 32'h3879c67b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f2; din <= 32'hb9ae00ca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c9; din <= 32'hc7dcdbf5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09c; din <= 32'h70d300e1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h366; din <= 32'h7e9822e3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a7; din <= 32'h907cb635;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28f; din <= 32'h050a4be0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a6; din <= 32'hc7d5ed2d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h333; din <= 32'hb6b7d4a7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h136; din <= 32'hce24795d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h256; din <= 32'had819db5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h099; din <= 32'h0917bb52;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h323; din <= 32'h57dc33bb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b4; din <= 32'h163f107b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25c; din <= 32'hfd334895;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b0; din <= 32'he8ffa3db;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3df; din <= 32'h2a57cdff;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a5; din <= 32'hf23cacba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h222; din <= 32'h8ee81e6c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00a; din <= 32'h2a617004;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31a; din <= 32'h33710bb3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h111; din <= 32'h3d0042cb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e8; din <= 32'ha029ef41;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h008; din <= 32'h05a5a320;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bf; din <= 32'hfedba3b3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h134; din <= 32'h2ecd38eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h206; din <= 32'h7f861e37;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h097; din <= 32'h2d5448f0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30a; din <= 32'he0d2be4f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ac; din <= 32'h787ccabe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27a; din <= 32'h49ff309a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h039; din <= 32'hd232dde0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ea; din <= 32'h8abb2085;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ea; din <= 32'h25eddf64;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26b; din <= 32'hb01c3dee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07c; din <= 32'h2bf29e53;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h370; din <= 32'h20096a91;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bd; din <= 32'hdf6974c3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e3; din <= 32'hf1b9b632;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02b; din <= 32'hd3887801;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h318; din <= 32'h0883fd72;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13d; din <= 32'hd6d0210e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c9; din <= 32'hcb81c4eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h060; din <= 32'hf30e1c47;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30d; din <= 32'h67d05889;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h181; din <= 32'h7c868c7b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f6; din <= 32'hc8b747c7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h098; din <= 32'h95d6a2c4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31a; din <= 32'h7f5ce43c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fd; din <= 32'h5ce2bbe3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e0; din <= 32'hc003b2a9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h019; din <= 32'hd39f3806;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h323; din <= 32'h477cfce1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ec; din <= 32'h81afdc48;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28c; din <= 32'h127ad4ad;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02c; din <= 32'hdda4968a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a9; din <= 32'h75b08d42;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c4; din <= 32'he24c7032;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21f; din <= 32'h3069e64b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05a; din <= 32'hdfbc6298;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h309; din <= 32'h3910ee3d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h199; din <= 32'hb6ef3494;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c9; din <= 32'hf6370890;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b3; din <= 32'hec00416d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ff; din <= 32'h31222e02;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14a; din <= 32'h4101f2c3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f5; din <= 32'h94075971;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h030; din <= 32'hd74f958b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33b; din <= 32'h42d956bb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h163; din <= 32'h0b165a4c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c0; din <= 32'h7518097e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01b; din <= 32'hf85886b9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35d; din <= 32'h9cad554f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bd; din <= 32'hd9838dc9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h215; din <= 32'hd57f4cc7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07b; din <= 32'hd2001dc0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h303; din <= 32'hd29781f3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cf; din <= 32'h33316397;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h225; din <= 32'h528bec95;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0dd; din <= 32'h1f9b2c50;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ba; din <= 32'hf0e5dfe5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ab; din <= 32'h0f4f6b21;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h233; din <= 32'h1bb9532c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h062; din <= 32'h9f56d5ad;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34c; din <= 32'he82712c4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h178; din <= 32'hbf682b7e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d0; din <= 32'hac451232;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b9; din <= 32'h19d746e4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32e; din <= 32'h47284431;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h190; din <= 32'ha616abf3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h287; din <= 32'h6d1f01d5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h012; din <= 32'h9c3f6a5f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39c; din <= 32'hade2af29;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h179; din <= 32'h14b88b79;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d1; din <= 32'h5e3b4c8b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h001; din <= 32'hd5ea6a08;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bf; din <= 32'hef754425;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h173; din <= 32'hc3712471;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29a; din <= 32'h9ebb0437;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c6; din <= 32'h0681fe02;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h365; din <= 32'h5bd958de;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fc; din <= 32'h9c4e92a3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b3; din <= 32'h7480ae53;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h059; din <= 32'h91ce45ec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h328; din <= 32'h2ce6c680;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h101; din <= 32'he8a3e30e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h204; din <= 32'hfff1053a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08e; din <= 32'hdfc811c8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e7; din <= 32'h45859b9e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bc; din <= 32'h0a333653;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h203; din <= 32'hed467b2f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h086; din <= 32'h508bab2a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cc; din <= 32'hee2787d5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h136; din <= 32'h0c19333d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f0; din <= 32'hb3817655;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h011; din <= 32'he18260c8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h311; din <= 32'hd1ecb665;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h118; din <= 32'hb4a26ba9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h212; din <= 32'hf5d92bfc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h089; din <= 32'h51c45e72;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3be; din <= 32'h0c4b0af3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c2; din <= 32'h418945eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h296; din <= 32'hb55bf103;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h004; din <= 32'ha21ae8bb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h396; din <= 32'h0ff643be;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h168; din <= 32'hc5859563;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24a; din <= 32'h300039f9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h091; din <= 32'h9c32d19b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30d; din <= 32'h0b72d103;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h145; din <= 32'h84b5cb89;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2da; din <= 32'h8101d0c2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h048; din <= 32'hbf2adb9d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30f; din <= 32'h5e25fa24;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1eb; din <= 32'h3d4218ec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27f; din <= 32'h160980f3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e5; din <= 32'haefa1dcf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37f; din <= 32'hfc6d0cd1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10a; din <= 32'ha25f1fd6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2af; din <= 32'h31a6b8fb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h001; din <= 32'h7980e758;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h351; din <= 32'hb84c9c99;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b8; din <= 32'h830ca135;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c3; din <= 32'h06de4ea6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08d; din <= 32'h53a5c5a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34e; din <= 32'h2d05eff0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h176; din <= 32'hdb005d40;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23a; din <= 32'h0e923a67;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h082; din <= 32'h30b8a54f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36e; din <= 32'h0459284c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19f; din <= 32'h0d84955d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ee; din <= 32'hc6fadab8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h086; din <= 32'hf605018e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c6; din <= 32'hcc573260;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h150; din <= 32'h2db01bf3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20d; din <= 32'h314e64cf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fa; din <= 32'hb5391b3c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ee; din <= 32'hba672a4f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a8; din <= 32'hf4aeac2e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h228; din <= 32'h30cd5d3f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h030; din <= 32'hb3ce832a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bd; din <= 32'h8c0c68e0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a1; din <= 32'h34ce6e01;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22f; din <= 32'h44acdf8b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a9; din <= 32'hf8eb5dea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cb; din <= 32'h5cb1dca8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16a; din <= 32'hc842ac07;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h288; din <= 32'h4da03532;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01f; din <= 32'h8f951aee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h353; din <= 32'h010e4ece;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h147; din <= 32'h38b0ac25;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b3; din <= 32'h1d92c462;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d1; din <= 32'hcdb81646;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36e; din <= 32'h415a0bdd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h145; din <= 32'hf7f5bc51;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20f; din <= 32'h3627b6eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h046; din <= 32'h28bbaac0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30c; din <= 32'hda2beb5f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h157; din <= 32'hefb68e31;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h225; din <= 32'h41fcac4e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d4; din <= 32'h29aa4a95;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b5; din <= 32'hc01d185e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h191; din <= 32'ha5563a8f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d4; din <= 32'hc56bdc95;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a8; din <= 32'h0653ab9e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b9; din <= 32'haffff32a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18e; din <= 32'hf4069a66;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f2; din <= 32'hc6ccbe6b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04f; din <= 32'h619dcb7a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h303; din <= 32'hf1eada21;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d8; din <= 32'h26541073;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b4; din <= 32'h1c9dfd6e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c8; din <= 32'he62e3293;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30a; din <= 32'h9215d40f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1dc; din <= 32'h02c8ce22;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27b; din <= 32'hc63f2b7b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08c; din <= 32'h9bb32ea6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37d; din <= 32'h23e33018;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h105; din <= 32'hba89f9f9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23e; din <= 32'h8e4b5990;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01d; din <= 32'h55cc25f4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3de; din <= 32'h31f37e3d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h186; din <= 32'ha661793f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c3; din <= 32'h272c6fdd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h082; din <= 32'h901582b4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32f; din <= 32'hea72e62a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h139; din <= 32'h7be96d4d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e8; din <= 32'h69ef438c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a6; din <= 32'hf2774a42;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a0; din <= 32'h8b4a246f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17a; din <= 32'h10712097;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ce; din <= 32'h7dd4ea6f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h009; din <= 32'ha1796122;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f5; din <= 32'h943cb90a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1aa; din <= 32'he83a215b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e3; din <= 32'h10638dde;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06e; din <= 32'h178be54e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a3; din <= 32'h7a8725b5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12c; din <= 32'h91178abe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24a; din <= 32'h3ac90471;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02e; din <= 32'hede01360;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35f; din <= 32'h1339412b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h169; din <= 32'h332f2aa5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24b; din <= 32'hdb0b8259;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f5; din <= 32'h05e31a4f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39d; din <= 32'h9af2538b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19b; din <= 32'hcb27c106;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h271; din <= 32'hc6b571d7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h041; din <= 32'ha25a8c92;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35a; din <= 32'hba9b6355;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c1; din <= 32'ha8f7678f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f6; din <= 32'h6dc32921;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h050; din <= 32'h6ad2ec1f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h317; din <= 32'h491c7b86;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h185; din <= 32'h0307887d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h261; din <= 32'hb53d00b2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b6; din <= 32'h90a1dca1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b6; din <= 32'h9122b13b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1be; din <= 32'h50d8bf2c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h256; din <= 32'hd55b7287;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h007; din <= 32'hc1329c86;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bb; din <= 32'h89e95298;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h161; din <= 32'hd19166ed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a8; din <= 32'h2250cb01;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h014; din <= 32'hb5b91004;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ed; din <= 32'hc9e172c6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cf; din <= 32'hab122b54;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h232; din <= 32'h4407e48e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f6; din <= 32'h9a773c7d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h357; din <= 32'h5d9e083f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f5; din <= 32'h5a5ceb95;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2af; din <= 32'h1f2ef071;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h097; din <= 32'h6c8a337a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h323; din <= 32'h89533e57;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b3; din <= 32'h2717dfb9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29c; din <= 32'h8ca6bcdf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01e; din <= 32'h91967655;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ac; din <= 32'hb37ae123;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13b; din <= 32'h202db89e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28c; din <= 32'h21867216;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0af; din <= 32'hfb0a9e44;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h397; din <= 32'h799f6f68;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h113; din <= 32'h97679eea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h239; din <= 32'h96f49b5b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a9; din <= 32'h977a119f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h363; din <= 32'h305565ed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h122; din <= 32'h07581ed5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e9; din <= 32'hcbe962d5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05c; din <= 32'h081c376f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h399; din <= 32'h10560129;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h156; din <= 32'hf642187c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a1; din <= 32'hb114c27a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h034; din <= 32'h3ce2113d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c4; din <= 32'h9b83f741;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1df; din <= 32'hde56885a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h201; din <= 32'hc53056b2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03e; din <= 32'haad8f2df;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34d; din <= 32'h319b9f94;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ae; din <= 32'hfd95bd28;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27c; din <= 32'hcea98016;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05d; din <= 32'h29e65b7a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30c; din <= 32'h68ff6397;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cc; din <= 32'h7813bbae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h269; din <= 32'h4226288d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h019; din <= 32'hec12e159;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e5; din <= 32'hcf051bb8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h124; din <= 32'h22a9772d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h210; din <= 32'he75142bf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01c; din <= 32'hd623cf44;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h371; din <= 32'h59e7625e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h175; din <= 32'ha2b9ccc7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d1; din <= 32'h240cf8d2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07f; din <= 32'hadd59ab4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bd; din <= 32'h4c2d591b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b4; din <= 32'h0e4dfc6d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h287; din <= 32'h3db85702;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f1; din <= 32'hb9bf87fa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h323; din <= 32'hd165b7ff;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ed; din <= 32'hf576bc3c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h291; din <= 32'h5ba36795;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h090; din <= 32'h583a8707;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bd; din <= 32'h5bf6cb07;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ff; din <= 32'hd6adb9d9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h253; din <= 32'hd1395157;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05b; din <= 32'h88471524;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e0; din <= 32'h550a2c77;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h118; din <= 32'he051ccf7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d3; din <= 32'h386d10be;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03b; din <= 32'had0c2dc6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cc; din <= 32'he1744afe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h183; din <= 32'h99b4c698;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e9; din <= 32'h8480f71d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h011; din <= 32'h052f761f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3eb; din <= 32'h7a707220;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h104; din <= 32'h70baf98d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e2; din <= 32'h44a76592;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h033; din <= 32'hb6b8f5f3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h374; din <= 32'h8698aaa1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10b; din <= 32'ha92d17b7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h270; din <= 32'h7671a781;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h050; din <= 32'heb0a64a2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34a; din <= 32'h1f2615e4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h140; din <= 32'h586e2491;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22c; din <= 32'h26782cb9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02f; din <= 32'ha4cf9a35;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h379; din <= 32'hf8e38fe1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ad; din <= 32'ha0e400be;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21c; din <= 32'hdc912043;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h081; din <= 32'h0dbfdb14;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h332; din <= 32'h96fcf812;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c1; din <= 32'hc3969645;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ff; din <= 32'h6bbc9659;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02c; din <= 32'h5fa93be4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e9; din <= 32'hc82a393e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h109; din <= 32'h86c78c9f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f2; din <= 32'h3cd5fb6f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00a; din <= 32'h795f9195;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31c; din <= 32'h29169e2f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1dc; din <= 32'hbdbffa94;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h297; din <= 32'hcf198d3b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h088; din <= 32'h0fd9d201;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a7; din <= 32'ha405f0e3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d2; din <= 32'h8c0c77c6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h290; din <= 32'h1147414d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02c; din <= 32'h935e4415;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h326; din <= 32'he4f42915;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e5; din <= 32'h4f18e98e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h259; din <= 32'hc3da27fc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ea; din <= 32'h49fc5dcc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h328; din <= 32'hb0e2090e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cf; din <= 32'h18a9ce8b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2dd; din <= 32'h6bc08e19;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cd; din <= 32'h4b1e4700;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37b; din <= 32'h66016564;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h191; din <= 32'h4cbe9b4c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h260; din <= 32'hc5b88e82;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f1; din <= 32'hb92b3a1e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35d; din <= 32'hfd53c095;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e6; din <= 32'hf518c044;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28f; din <= 32'hc72ab023;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e6; din <= 32'h34e66d96;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h313; din <= 32'h09a3d9a5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18f; din <= 32'h3f1fc499;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c1; din <= 32'he0aa7425;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01d; din <= 32'h51306e7d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cb; din <= 32'h6ed878fc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ea; din <= 32'h91d3dc13;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21f; din <= 32'h564c0e2a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09d; din <= 32'h799c1384;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h366; din <= 32'h5c81d940;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bd; din <= 32'h8bf77ddc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h203; din <= 32'h9fd454f5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h050; din <= 32'h9efb0ab1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f2; din <= 32'h2a236280;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18b; din <= 32'hd9dee40c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c1; din <= 32'ha3f3cce3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04c; din <= 32'h6b5b01a3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33d; din <= 32'h5a163e99;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h121; din <= 32'hdc8ddd16;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ac; din <= 32'h6a205579;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00a; din <= 32'h61c96966;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ab; din <= 32'hd855c170;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12c; din <= 32'hfd27a8a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2de; din <= 32'hcaa0e3bc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b3; din <= 32'he674ce7f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h371; din <= 32'h2ce1226a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h197; din <= 32'hb8da1219;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25c; din <= 32'h1460c839;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h048; din <= 32'h98aec5e3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h341; din <= 32'he926e741;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c4; din <= 32'h416ac11a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bf; din <= 32'haa416ad9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h070; din <= 32'h8e9f8ce1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c0; din <= 32'hea456d97;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h198; din <= 32'h02ee0461;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h207; din <= 32'hf597bd3c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h017; din <= 32'he3774940;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b2; din <= 32'h6258607e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h133; din <= 32'h579bf2d7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26d; din <= 32'h10bd90c6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c2; din <= 32'hcf28667e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f1; din <= 32'h70f5c333;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18f; din <= 32'h4ea8d34a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h251; din <= 32'h77f95dd7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05b; din <= 32'h737e605d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34d; din <= 32'h7ae59eaa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18d; din <= 32'h9b716606;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h212; din <= 32'hfe7e815e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ad; din <= 32'hba6dd257;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34f; din <= 32'hf291da9e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17c; din <= 32'h4bcce4d4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h214; din <= 32'hb2fe72de;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ef; din <= 32'hefaa43d9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h389; din <= 32'hf1626435;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h198; din <= 32'h29535555;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29a; din <= 32'h8cdee8ac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a5; din <= 32'h5ef9459f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39b; din <= 32'h9f23097f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h164; din <= 32'hb540c045;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h238; din <= 32'hdd5f2b80;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ae; din <= 32'h6567d4e6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d5; din <= 32'haf2e847a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13d; din <= 32'hc5de0488;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h228; din <= 32'h54a25ecf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h052; din <= 32'hb7a1d0b2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30e; din <= 32'h1a0fa951;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h182; din <= 32'h246ae89e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21d; din <= 32'ha5cc3ee6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f5; din <= 32'h78511132;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31d; din <= 32'h9599801c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h106; din <= 32'hd73ffdeb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h270; din <= 32'h53d59ccd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cb; din <= 32'hdc2795b1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ba; din <= 32'h14c40444;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ab; din <= 32'hd730d793;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h272; din <= 32'h34b88ba6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02a; din <= 32'h0889e62b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ec; din <= 32'ha9232b5c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h115; din <= 32'h864469bc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d5; din <= 32'h3de6911f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h023; din <= 32'hf4acffc5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e4; din <= 32'h8f4cb94a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a8; din <= 32'h5d823730;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h242; din <= 32'h3cc0851e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0db; din <= 32'h61ad0719;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32a; din <= 32'hb7bed95a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b4; din <= 32'h18cd9ede;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d8; din <= 32'h44cd6b67;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f3; din <= 32'h04bcd5d4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h385; din <= 32'h4842e86f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d7; din <= 32'h57d5b13d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22a; din <= 32'h2f2d1243;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c2; din <= 32'hdcd02fc8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b0; din <= 32'h96ec9b5c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b9; din <= 32'h9ed3b075;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h285; din <= 32'h2e4b6c32;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h085; din <= 32'haf12f872;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h341; din <= 32'h52e756a1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h120; din <= 32'h1f95bfed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h204; din <= 32'h0a765ead;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02a; din <= 32'hfc309898;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h399; din <= 32'h445120fd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c4; din <= 32'h6398b2b2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h285; din <= 32'hd0a7d34d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f4; din <= 32'h1f52122a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33c; din <= 32'h2e548ebf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h127; din <= 32'hf630979f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h244; din <= 32'h63302a9a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06b; din <= 32'h0acc607d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39a; din <= 32'h61e05811;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c6; din <= 32'ha7caef1d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20f; din <= 32'h269bc0ed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d4; din <= 32'h43f5e095;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h335; din <= 32'hfbf1b50c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a4; din <= 32'h9825f825;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h293; din <= 32'hf5892ac0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h058; din <= 32'hc5edd9c6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37f; din <= 32'h16483c2a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fe; din <= 32'h71178a40;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h215; din <= 32'habffc0b6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05b; din <= 32'h35cad7f7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h302; din <= 32'h9cf80ffd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h115; din <= 32'he5c0eb77;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h234; din <= 32'h2d645f0a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h044; din <= 32'h84901551;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39b; din <= 32'hb97d0d05;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bc; din <= 32'hb62b62d3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h207; din <= 32'h752aaa26;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04f; din <= 32'h6b06ba90;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h335; din <= 32'haee62241;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e0; din <= 32'hed8b0427;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e6; din <= 32'h522e1c01;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h055; din <= 32'heeb8ee55;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f5; din <= 32'hd7af2bc9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c9; din <= 32'h4a5b0778;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h275; din <= 32'h420b3a4c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0de; din <= 32'ha9ef9190;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h324; din <= 32'hf8740bc8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1dc; din <= 32'h173ce5e8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21a; din <= 32'h4ca5b5bf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h073; din <= 32'h6fc0cce5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31c; din <= 32'h527bbd16;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15e; din <= 32'h961b4b72;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27a; din <= 32'hf89b03c0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h011; din <= 32'hc633edd8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fc; din <= 32'h503a1af6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17c; din <= 32'h0243e18c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d8; din <= 32'h6729574e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09e; din <= 32'h398eb5d3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31e; din <= 32'h906ce673;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16a; din <= 32'h082b8bc5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c6; din <= 32'hdf7b5ed2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d4; din <= 32'hf7b52ec5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h341; din <= 32'hff7af22c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h131; din <= 32'h337b7028;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f2; din <= 32'h92dd04d2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05e; din <= 32'hf08aa87c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h319; din <= 32'h9634e86e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1af; din <= 32'h17dd29be;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28b; din <= 32'hcadb7f5b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h081; din <= 32'h17078309;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fa; din <= 32'hc8571985;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16d; din <= 32'hd99d31ae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24a; din <= 32'hca7b32c5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h098; din <= 32'h9695c4e6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h335; din <= 32'hf06c0329;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12f; din <= 32'hca00f7b4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h240; din <= 32'h323e7f1e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bf; din <= 32'h1570e13a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b1; din <= 32'hc19d4f02;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h134; din <= 32'hed258634;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e1; din <= 32'h1044d03b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h051; din <= 32'hb8075381;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h328; din <= 32'h92c76267;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bc; din <= 32'h8af2e43e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h255; din <= 32'h7d6d0dcf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cb; din <= 32'h7a514a68;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h360; din <= 32'h36cf0ae4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17f; din <= 32'h947bf3ce;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23b; din <= 32'h1112dd4d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h007; din <= 32'hef8b27a8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d0; din <= 32'hef51fa32;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h143; din <= 32'he0fbb11a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c9; din <= 32'h11f4eb47;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ab; din <= 32'hd3b10c29;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cb; din <= 32'h4725eca2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17e; din <= 32'haaedb220;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h261; din <= 32'h297dd431;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h093; din <= 32'hb9df201c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d4; din <= 32'hbfbce258;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cf; din <= 32'h2a31ce70;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20d; din <= 32'h00feb308;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03b; din <= 32'hfe0bee1e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bb; din <= 32'hc34a5eb7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17a; din <= 32'ha4a12ded;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h201; din <= 32'hd4b3a8f1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h081; din <= 32'h72e1b780;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3eb; din <= 32'h484bbd38;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cb; din <= 32'h1b7a7618;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h234; din <= 32'h9772eb09;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e7; din <= 32'he9549a29;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30d; din <= 32'hb9913c6c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h123; din <= 32'h5cfa4563;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26c; din <= 32'h1a2026ae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h066; din <= 32'h59b0574e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f3; din <= 32'h1e8cbc30;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18c; din <= 32'he8b2e926;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h292; din <= 32'h65f241a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h021; din <= 32'h8668d63a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ad; din <= 32'h7b50b5fa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h179; din <= 32'h7d8e4955;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28f; din <= 32'h2a3b4d8b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h061; din <= 32'h3786bebd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h398; din <= 32'h40da752b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h114; din <= 32'h5ac5b788;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29c; din <= 32'hb55f678f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01b; din <= 32'h51fad7d0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h386; din <= 32'h09a3d465;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15c; din <= 32'h045002bb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e4; din <= 32'h41563a94;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h023; din <= 32'h60dac9e5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ff; din <= 32'hf9babb6b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e1; din <= 32'hcd923dc8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2be; din <= 32'h55d13cfd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h027; din <= 32'h5e0c2221;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3df; din <= 32'he9595e99;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19d; din <= 32'h43be0ab4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h299; din <= 32'he6d72f4e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e3; din <= 32'hfa16a868;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3af; din <= 32'h919524a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19d; din <= 32'hbd90fcf2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22b; din <= 32'h5c826cc6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09c; din <= 32'h45658b91;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fd; din <= 32'h4e9b17da;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bc; din <= 32'h73b44983;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21e; din <= 32'h820fcb3b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08b; din <= 32'h11d37612;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e9; din <= 32'ha9128ae6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18f; din <= 32'h77322027;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h218; din <= 32'habaf4a32;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c2; din <= 32'h52b36140;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34f; din <= 32'h64ab765a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h110; din <= 32'he0ca71a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h269; din <= 32'h228b80a4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d3; din <= 32'hf8445988;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h352; din <= 32'he2938e4c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13f; din <= 32'h08bbfb13;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h247; din <= 32'h002bc67a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fc; din <= 32'h4c35e39e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b8; din <= 32'h8958ee89;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ad; din <= 32'h50d4faec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b3; din <= 32'h80ef664f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f3; din <= 32'hdb76400d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e5; din <= 32'he1f64638;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d6; din <= 32'h0f8c1d1c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2eb; din <= 32'h9a3e5495;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f2; din <= 32'h43257110;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ff; din <= 32'h753c14b6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13c; din <= 32'he0116af5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h292; din <= 32'h16a23ce6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e5; din <= 32'h800ab4ff;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h371; din <= 32'h2aace610;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b8; din <= 32'h84f85cb9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h251; din <= 32'h0d2cd311;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06f; din <= 32'h1edcccb2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f6; din <= 32'h12da4600;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h177; din <= 32'h9813d2c3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h256; din <= 32'hd8dd3fae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h041; din <= 32'he3ea366e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34e; din <= 32'h8702dcf6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f1; din <= 32'h49496c12;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h294; din <= 32'h7955d370;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e9; din <= 32'h69cf65ed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h335; din <= 32'h324a3837;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12f; din <= 32'h61e538d3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h289; din <= 32'h212043df;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03e; din <= 32'hb9e84193;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3eb; din <= 32'hcbc9aef0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h187; din <= 32'hc06b1c49;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25d; din <= 32'hc9592cbc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09a; din <= 32'h75da1336;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3db; din <= 32'h7956784e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18c; din <= 32'h5d8de125;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h260; din <= 32'h62288a54;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e1; din <= 32'h2bd0b520;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d6; din <= 32'h39766f39;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h132; din <= 32'h796cccc6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h244; din <= 32'h1df19491;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h086; din <= 32'he00b14c4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h383; din <= 32'hfec796c3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h129; din <= 32'hb4bb7783;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h264; din <= 32'h9e1dff09;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a9; din <= 32'h795d6131;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c4; din <= 32'h6a61ed23;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d8; din <= 32'ha9352b3a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h215; din <= 32'h477532bf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h026; din <= 32'h6451e80b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h337; din <= 32'h9c7365f1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10f; din <= 32'h90aace69;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cc; din <= 32'h1ed98da4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h032; din <= 32'hbc77f948;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a9; din <= 32'h753bb348;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fb; din <= 32'hc331029d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24b; din <= 32'h8236ad71;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cd; din <= 32'hc362aa4d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35e; din <= 32'hc61e8fa8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b2; din <= 32'h2430ce17;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h221; din <= 32'haab120f8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a9; din <= 32'hd9b4d788;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30e; din <= 32'hacfba0d7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c9; din <= 32'hacc7a143;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cc; din <= 32'he0c3fcee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05d; din <= 32'h72545706;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h307; din <= 32'hb089b1da;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h162; din <= 32'he3cf4849;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h206; din <= 32'h9b97eebb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h011; din <= 32'h4b6852f3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31e; din <= 32'h85cf4927;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h169; din <= 32'h9adae400;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h216; din <= 32'hf6e4c0d9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08e; din <= 32'h6b6a759a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h388; din <= 32'hf1c1c478;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14b; din <= 32'h079bd67b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e2; din <= 32'h125e3af5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h009; din <= 32'h6f6c1a27;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h391; din <= 32'h74ca34d7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h132; din <= 32'h03c5fbf8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h277; din <= 32'hd9fe30dc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03d; din <= 32'hf781f3f0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h348; din <= 32'h4ad08a96;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f5; din <= 32'hba5b3339;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h278; din <= 32'h5e313bf2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c4; din <= 32'he9ef381a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h336; din <= 32'he31c13a5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13f; din <= 32'he06a8b5d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h226; din <= 32'h3997bb05;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06e; din <= 32'hd6fadde8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ab; din <= 32'he3e8209c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h153; din <= 32'he009f7f6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h270; din <= 32'h2ffd0d7f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03f; din <= 32'h538b4081;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a4; din <= 32'h68a9b9de;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e0; din <= 32'hc7361379;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22d; din <= 32'he4bcfbae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h085; din <= 32'h3209de83;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39c; din <= 32'h70cc97b1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h128; din <= 32'he91ed0c7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h239; din <= 32'h8834c398;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h040; din <= 32'habed0b65;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bf; din <= 32'h6f5f2889;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16a; din <= 32'h8264dca3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b1; din <= 32'h1be8654c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03f; din <= 32'hadc9d2eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h356; din <= 32'h5ce6f639;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e4; din <= 32'h931830f1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22a; din <= 32'h65501f13;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02f; din <= 32'hc76c6e29;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h385; din <= 32'hd5b04a48;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f1; din <= 32'he2798a5d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h231; din <= 32'h3368491a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h062; din <= 32'h123c824c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fc; din <= 32'ha3a1c49a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ba; din <= 32'h2dc55fe9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h291; din <= 32'h625ad6d8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05c; din <= 32'h08bdc3a8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d0; din <= 32'h60811e4f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h171; din <= 32'h6c28dbb5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a8; din <= 32'h652809a7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c5; din <= 32'h1c1c4c2c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h322; din <= 32'hb42058f4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18f; din <= 32'hc6624a6b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c9; din <= 32'h4e0ad180;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01e; din <= 32'h08c69f4e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d1; din <= 32'ha10f224a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h176; din <= 32'h96b3fbcf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b0; din <= 32'h5d79f4ee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h025; din <= 32'hf51b63a1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39d; din <= 32'h09a39354;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c9; din <= 32'hc7ba8518;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h259; din <= 32'ha2e870f7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09f; din <= 32'hc79d1224;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cd; din <= 32'ha2f67566;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h176; din <= 32'h52aac04f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f2; din <= 32'hc49373d8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h062; din <= 32'h1015d613;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34d; din <= 32'h1c0d978d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h103; din <= 32'he3a900cb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h200; din <= 32'hd5ead677;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h030; din <= 32'hb3451415;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h300; din <= 32'ha74cf668;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h196; din <= 32'h4472d6f8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h257; din <= 32'hf77f3e4a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07c; din <= 32'h81898865;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d0; din <= 32'h10d69713;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h168; din <= 32'hd5476957;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ac; din <= 32'h7d223d58;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07c; din <= 32'hf58e28bc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34b; din <= 32'hb787eda3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fb; din <= 32'ha60500ac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a3; din <= 32'h5e0719c4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b7; din <= 32'h6f641f6d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35c; din <= 32'hff594f42;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h178; din <= 32'hb44da34e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h258; din <= 32'h7b15f8d3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d7; din <= 32'he1575f09;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h341; din <= 32'he66679c6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10c; din <= 32'he84fa5a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ba; din <= 32'h1b91e6be;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h019; din <= 32'h6aa1de2e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35d; din <= 32'hbb5f8f2b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cd; din <= 32'ha81c12c4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h277; din <= 32'hbe20f3eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04b; din <= 32'h0e9d713f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c2; din <= 32'h654ae83a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h173; din <= 32'h02b630cf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b1; din <= 32'h2dec6bf6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h070; din <= 32'h0950d3a9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cb; din <= 32'h050955e1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13a; din <= 32'h0620aeab;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c6; din <= 32'haec191d7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h026; din <= 32'ha9ea2776;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ab; din <= 32'h137a9a0d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h123; din <= 32'hdb1bc91b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h217; din <= 32'h67b66809;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h055; din <= 32'ha1a35d3d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39d; din <= 32'h01cd94d2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e4; din <= 32'h18b3e682;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20c; din <= 32'h1c362211;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h054; din <= 32'h7a5666f6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h309; din <= 32'h105caa8e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b3; din <= 32'h3d9b2f1d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h244; din <= 32'hd4facd4a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h055; din <= 32'hbd4b91b0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h379; din <= 32'h91b66ad5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h110; din <= 32'h721eb3d6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h261; din <= 32'hb44bd8fc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0eb; din <= 32'h425dc078;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h364; din <= 32'h37cfc2bf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15a; din <= 32'h88dff6f7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28c; din <= 32'hf1b25418;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e5; din <= 32'ha6b3f874;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32f; din <= 32'h9ad8cbb8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19b; din <= 32'hf94e7964;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23e; din <= 32'h4c7937ca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h086; din <= 32'hdba4fe05;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31f; din <= 32'ha0f455ac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h121; din <= 32'h5e64f514;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a7; din <= 32'haae3dc86;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e9; din <= 32'had554263;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h311; din <= 32'h23b2d671;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12d; din <= 32'hf7b2e166;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h226; din <= 32'ha5e07830;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c3; din <= 32'hc880b676;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f0; din <= 32'h7e88b454;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d2; din <= 32'h5da1b410;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20b; din <= 32'h37e8a163;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06a; din <= 32'he15c080e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ed; din <= 32'hd97e7209;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fa; din <= 32'h4d0ac817;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a9; din <= 32'hc81469aa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03e; din <= 32'h036bf55b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h354; din <= 32'h9596e940;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h171; din <= 32'hc9f16fa4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2dd; din <= 32'he556e830;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04a; din <= 32'h391f3e5d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33f; din <= 32'h2945b508;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17b; din <= 32'h24e2db2c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h258; din <= 32'hd06a946c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h024; din <= 32'h999c018c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31e; din <= 32'h31632028;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h176; din <= 32'h8e53c147;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23d; din <= 32'h28d93a05;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h087; din <= 32'h68789dd6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3be; din <= 32'h1fdc4003;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b9; din <= 32'h2cd3f851;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ba; din <= 32'h59a67932;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ab; din <= 32'hec099d5d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h332; din <= 32'h31d51b33;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f0; din <= 32'h2962cdf9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h239; din <= 32'h5cc056e1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c9; din <= 32'h58b1c1c9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34d; din <= 32'h0b160db9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1df; din <= 32'h37b2ee04;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h293; din <= 32'hf8e64df5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ad; din <= 32'h2bc035fa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33d; din <= 32'h5ebc5a1c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12d; din <= 32'h0e49dc26;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25a; din <= 32'h46f24a82;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h081; din <= 32'h475daf30;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d6; din <= 32'h7aaec978;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h112; din <= 32'h960b4477;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h225; din <= 32'h06626080;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08e; din <= 32'h87051eac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30b; din <= 32'h7ce4b164;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h158; din <= 32'hc112e9c9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h262; din <= 32'hc008a41f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c9; din <= 32'h696b2127;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c3; din <= 32'h59a56026;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14c; din <= 32'h4a6fdb8e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a1; din <= 32'hf65e90e5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d2; din <= 32'h5e41c5bf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cb; din <= 32'h6c9dc7ac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ea; din <= 32'h0225534e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25f; din <= 32'h1d7a43dd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h025; din <= 32'h43755a34;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33b; din <= 32'h1a921287;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fd; din <= 32'hcdb03044;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h212; din <= 32'ha3fb0ae2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h076; din <= 32'h4d2602ac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h363; din <= 32'h5859364d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fb; din <= 32'h0f99ec96;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h299; din <= 32'h8bc1aad4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01e; din <= 32'h5f00c2c5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h368; din <= 32'h99a11c6d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h184; din <= 32'he7ea6fe1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c2; din <= 32'h5b462e20;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ab; din <= 32'h264f3ab7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f9; din <= 32'ha7e2ac34;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h175; din <= 32'hc975bd69;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h226; din <= 32'h808e6cce;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fb; din <= 32'hdeede0fe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h380; din <= 32'h7ade6f47;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h192; din <= 32'hfb236cfa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h239; din <= 32'h9a1ae6d2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d9; din <= 32'h335ad673;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h353; din <= 32'h6a1af1de;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19a; din <= 32'hf078e0a1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ea; din <= 32'hdf52e92f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h057; din <= 32'hea00ce56;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d2; din <= 32'h9c829a58;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h168; din <= 32'h477687cb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e8; din <= 32'hcd4630dd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h092; din <= 32'hd4b86fa3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ce; din <= 32'h0f55cada;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15f; din <= 32'hd58a9f83;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h217; din <= 32'hc6f4db83;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h085; din <= 32'hb854a313;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h336; din <= 32'hd5b6d043;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h124; din <= 32'hd88602c8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24e; din <= 32'h36dd11f4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h037; din <= 32'h475201de;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30f; din <= 32'h73f90821;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1de; din <= 32'h07e7f047;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22a; din <= 32'h5f4008f1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h051; din <= 32'h6b77e6b6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ca; din <= 32'hb36b3f4b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13c; din <= 32'h17228982;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e3; din <= 32'ha27ad6c4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b3; din <= 32'he634e53d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h386; din <= 32'h84bb783e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h124; din <= 32'hbcced8b1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29a; din <= 32'h9c9964f2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h030; din <= 32'h46f1d205;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h350; din <= 32'h59c6000b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h162; din <= 32'he1d86743;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23b; din <= 32'hcb0e214f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h094; din <= 32'h559bd4ea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h325; din <= 32'h0eedbe06;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a9; din <= 32'h4774844e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c0; din <= 32'hae96f813;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h053; din <= 32'h2503ebc2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h318; din <= 32'h9fb3cafa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cc; din <= 32'h2767d973;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2de; din <= 32'hb8e449c7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06e; din <= 32'h7b92b2db;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e2; din <= 32'h5e937add;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19c; din <= 32'h3ddabb30;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2fe; din <= 32'h46d4d845;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04b; din <= 32'h9ff43f5e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e2; din <= 32'hb6dc0f8c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h142; din <= 32'h05f592d8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ad; din <= 32'h353de0d8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c8; din <= 32'hd7455db6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h353; din <= 32'h60ddde28;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12b; din <= 32'h35ed7e1a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h290; din <= 32'h6a52ede2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03e; din <= 32'h958db32f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37b; din <= 32'h7745c344;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11e; din <= 32'h1a25d45a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21b; din <= 32'h6e71386d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0aa; din <= 32'hbe9383ef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h334; din <= 32'h6181545b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cb; din <= 32'ha2e075b1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h261; din <= 32'hdc6d190a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h061; din <= 32'hfb65ed4b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e8; din <= 32'h6cf967af;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h181; din <= 32'hfe79addf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bf; din <= 32'h613696e8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h086; din <= 32'hdea6643a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h349; din <= 32'h5cce8a5a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a6; din <= 32'h0a195f51;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h286; din <= 32'h60b2b37f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ad; din <= 32'hbb2731c2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b1; din <= 32'h279156af;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h109; din <= 32'h2bd0fd4a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24c; din <= 32'hebe32777;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d7; din <= 32'h5fc813af;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b5; din <= 32'h23d2b288;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a5; din <= 32'hf39460b4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bf; din <= 32'h0264bc47;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02d; din <= 32'h316399a8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h333; din <= 32'h2e956a13;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h198; din <= 32'h07ffcd76;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2eb; din <= 32'h811316c6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h038; din <= 32'h62afeb9e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h394; din <= 32'h9fe9182e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ea; din <= 32'h2254fac0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h240; din <= 32'hbc2dd1a4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00e; din <= 32'h5cab1af8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h382; din <= 32'h85cb376e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h123; din <= 32'h1108ec2f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h243; din <= 32'hd9ca1ee7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a2; din <= 32'h43c66706;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32b; din <= 32'hbca1e7c0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16d; din <= 32'h8a8eab7f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h204; din <= 32'hd294c2f1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d9; din <= 32'ha1163e92;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h356; din <= 32'hccb39acf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12f; din <= 32'hb89c50a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29f; din <= 32'h566c0eee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h060; din <= 32'h0460c7ba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h322; din <= 32'hdf31174e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h184; din <= 32'hc2076ab9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f7; din <= 32'h46834e0e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d7; din <= 32'h5507544f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h303; din <= 32'h8e3bb7c7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1da; din <= 32'h89fc499c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b1; din <= 32'h4504f8f1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09d; din <= 32'he071d2d4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h388; din <= 32'he6c1f13c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h150; din <= 32'ha0c2cdcd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2be; din <= 32'h22aa5d6d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04b; din <= 32'h023ac0b7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31c; din <= 32'h4c3dc326;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h116; din <= 32'h79600e1d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ea; din <= 32'ha354ddd8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b6; din <= 32'hfbe99b27;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h335; din <= 32'hcc03cad2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17e; din <= 32'h000acdec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a1; din <= 32'hafc83b0c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h034; din <= 32'h72d3e197;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h379; din <= 32'h2bb85c72;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ee; din <= 32'h7296d66b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bd; din <= 32'h01af23b8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08c; din <= 32'h76d8779f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3dd; din <= 32'h963a4337;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h104; din <= 32'ha634fef0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h266; din <= 32'hc77b1731;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05e; din <= 32'h6466d608;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h311; din <= 32'h26ef6bcd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c5; din <= 32'h15d5ea6a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h289; din <= 32'hecedd664;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05b; din <= 32'h12e5356f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h313; din <= 32'hdbaf331e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e9; din <= 32'h70d12dea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20b; din <= 32'ha0b06f02;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c4; din <= 32'h1427a8ba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h302; din <= 32'h30476aa2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b7; din <= 32'hbcff33c6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h214; din <= 32'h5578d69b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bb; din <= 32'h83963e94;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h358; din <= 32'he77922fb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e3; din <= 32'h14ca9cdb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20d; din <= 32'h280f04c8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h045; din <= 32'hdc89f704;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36a; din <= 32'h26a0b9fe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h131; din <= 32'h2896cee7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h230; din <= 32'hbd520944;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d1; din <= 32'hc005dfe0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h373; din <= 32'h8e45ce7d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19e; din <= 32'h47b600a1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d4; din <= 32'ha03f375b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h055; din <= 32'h81d9a9bd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fa; din <= 32'hd628837c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14c; din <= 32'hf9a75ade;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c5; din <= 32'h6778a1f6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h007; din <= 32'hf74c1e30;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h322; din <= 32'hdbfa0173;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h180; din <= 32'h3c3fa195;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22a; din <= 32'h673b8a5d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h079; din <= 32'h48e9baba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cb; din <= 32'h293116b8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h141; din <= 32'h57ad2cfe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e3; din <= 32'h6dc5a3ee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e8; din <= 32'h84a2e42d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33b; din <= 32'h22069062;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h180; din <= 32'h1c809caf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h212; din <= 32'h8605f8a4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ba; din <= 32'hdbb503df;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ec; din <= 32'h14dcaede;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h156; din <= 32'h5bbf967e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ef; din <= 32'hfb8af153;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h068; din <= 32'h614fbc16;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c4; din <= 32'hb031a2ce;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b8; din <= 32'h89d4bd3f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h229; din <= 32'ha301d860;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h089; din <= 32'hfee1b473;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h334; din <= 32'hb67b28bd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18b; din <= 32'hf272af8e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2eb; din <= 32'h3a7952b5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02b; din <= 32'h3567f8cc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35e; din <= 32'h316c1e79;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a4; din <= 32'h3d962857;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20d; din <= 32'h00cd8e08;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c8; din <= 32'h802af6a1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fc; din <= 32'h0454d8e4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d6; din <= 32'h1cdb7f01;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h269; din <= 32'h19b21ce8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cc; din <= 32'h404b44e4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3de; din <= 32'h84fa3679;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h161; din <= 32'h894114f6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b2; din <= 32'h317522c2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h024; din <= 32'h5e82a2ac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h343; din <= 32'hf59789ba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15d; din <= 32'h22962005;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h219; din <= 32'hf0477903;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c5; din <= 32'h787fab53;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35b; din <= 32'h051e856c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13d; din <= 32'h07dd26f9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h254; din <= 32'h505c8e3a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05e; din <= 32'hcac6980f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h384; din <= 32'hdfeb801c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ce; din <= 32'h635a1d2c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h296; din <= 32'hb170762d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bb; din <= 32'h462da06e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a4; din <= 32'h519c7767;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d0; din <= 32'hc117e49b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bf; din <= 32'hc8060579;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01f; din <= 32'h942aa255;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h313; din <= 32'h3a5997db;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h144; din <= 32'h995fd80a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cf; din <= 32'h9b602613;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d8; din <= 32'h6b7e1b1c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h365; din <= 32'hd83c2fa7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ce; din <= 32'h88ddd14d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e5; din <= 32'h68ecf9c8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h032; din <= 32'h1273b1c3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h336; din <= 32'hac5321c5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h175; din <= 32'h0c162c0b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d0; din <= 32'h8a2f69c3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h022; din <= 32'h714dc325;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e7; din <= 32'h770fd77e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h182; din <= 32'he879f5da;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h270; din <= 32'hb06c6d3f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h021; din <= 32'h68388b82;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39f; din <= 32'hd75b40cf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17e; din <= 32'h7f392cb0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28b; din <= 32'h34aa8a10;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02f; din <= 32'h88040e85;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b5; din <= 32'h2787b1a7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h122; din <= 32'hfdbee01e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24d; din <= 32'hafcbae66;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h046; din <= 32'h26863378;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h331; din <= 32'hf19203b1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h157; din <= 32'h01b329c1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d0; din <= 32'h81d042bb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h057; din <= 32'h6992597d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h359; din <= 32'hbe877fdc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11f; din <= 32'ha7b8e3a4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e2; din <= 32'h92e03270;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fc; din <= 32'hefc343ef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d7; din <= 32'hd9c18127;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d1; din <= 32'h9df52767;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h210; din <= 32'heabf57eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h032; din <= 32'hb50baef6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cf; din <= 32'h84ae6028;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ad; din <= 32'hde5290e7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26a; din <= 32'h16f29e74;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e8; din <= 32'h1348339d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ac; din <= 32'h8e9e68f1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d4; din <= 32'h4b7a0aa4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h281; din <= 32'hd995ac93;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06b; din <= 32'hd6c7105f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h308; din <= 32'h2782ded4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h191; din <= 32'hec26db6e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24f; din <= 32'haacdba18;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h008; din <= 32'h7aedcc83;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34e; din <= 32'h18be8a5c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h141; din <= 32'h0c4cbc02;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20a; din <= 32'hbbe63482;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h020; din <= 32'h926cd40f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h350; din <= 32'h8be1804b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19e; din <= 32'h3a7e60f7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h211; din <= 32'h5dca3e57;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02b; din <= 32'h4a30489d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h312; din <= 32'hc968afa4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a3; din <= 32'h9317ebf3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2de; din <= 32'he564199d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h080; din <= 32'hf5997f92;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a9; din <= 32'h4cd816f6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17c; din <= 32'h5a31cd59;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22e; din <= 32'h6cf03564;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06b; din <= 32'hcb70058f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h308; din <= 32'h6b4757e4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10f; din <= 32'hedb2ffa3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h296; din <= 32'hb5f5aa7a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c3; din <= 32'hf4f62b07;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f3; din <= 32'h2ba5386f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11c; din <= 32'h7ce07ef1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24b; din <= 32'hb17cdaee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f4; din <= 32'hcc913e94;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d2; din <= 32'h5036f748;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10b; din <= 32'h64bc1f0f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20c; din <= 32'h80fd48f4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06d; din <= 32'hc728d8e8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h316; din <= 32'h984d8d8e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h176; din <= 32'h91326c9d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2db; din <= 32'h6b1e7f4f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h070; din <= 32'h7c6ae9be;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h359; din <= 32'haa2c35df;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10f; din <= 32'h2ba81f45;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h293; din <= 32'hbdc7f1fa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h021; din <= 32'h78b7a2fb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3aa; din <= 32'h01bd6070;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ac; din <= 32'hf2df6dd6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e3; din <= 32'h4a234c26;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04a; din <= 32'h7ba50947;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31a; din <= 32'hedb67991;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h159; din <= 32'hac32b45b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2fd; din <= 32'hef281e39;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h049; din <= 32'h43181818;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c1; din <= 32'h3024f816;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h111; din <= 32'h7c0e404e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c2; din <= 32'h83ea801d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h050; din <= 32'hdf178e85;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h387; din <= 32'hf63c9e43;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h129; din <= 32'h789a0964;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b9; din <= 32'hd79d3f7a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d5; din <= 32'he8e1cb43;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h314; din <= 32'h9c109cb6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h148; din <= 32'h463ee873;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20e; din <= 32'hb85ecf66;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02e; din <= 32'hc50bc245;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h328; din <= 32'hde9d75fd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13d; din <= 32'h8dd44232;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d5; din <= 32'hdcfd7717;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03b; din <= 32'h27f1d54c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h345; din <= 32'h509700e4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fa; din <= 32'h2ea1244e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e5; din <= 32'hd3843f01;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h087; din <= 32'h6a33e36e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h361; din <= 32'ha5c9442a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h168; din <= 32'he5b42c3d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h200; din <= 32'hfd54297f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cb; din <= 32'h7557c183;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h353; din <= 32'h31aecdb9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h127; din <= 32'h8cb52797;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bc; din <= 32'h9155e0df;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h079; din <= 32'h8ba1defc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h335; din <= 32'h8d443ae7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e3; din <= 32'hff3c99fe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25a; din <= 32'h36a43597;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h018; din <= 32'ha88801d5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d6; din <= 32'he18dba59;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e4; din <= 32'h247c48e2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d7; din <= 32'h176def25;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h047; din <= 32'h85c1031d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h388; din <= 32'hf7513a97;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13a; din <= 32'hc8a6fc53;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h256; din <= 32'hb4160fd2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a3; din <= 32'h5e6b55e7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33b; din <= 32'h21681c38;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1be; din <= 32'h85891b6f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h292; din <= 32'hfc13280e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h027; din <= 32'h088e4069;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ea; din <= 32'h76c061b3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h186; din <= 32'h7923d6dc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h285; din <= 32'h17a258db;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03d; din <= 32'hb7629b30;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h325; din <= 32'h51ec1e36;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12d; din <= 32'h3f25222b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h295; din <= 32'h4470626f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f1; din <= 32'h272c4faf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c5; din <= 32'h61eaf8b1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h143; din <= 32'h19d5d4d6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h274; din <= 32'h59b4d837;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e3; din <= 32'hb7a44291;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h303; din <= 32'ha806a19c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16e; din <= 32'hb5f0300e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d7; din <= 32'hb0cc72a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c9; din <= 32'h55db7d9b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d2; din <= 32'h4a735481;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17a; din <= 32'h60bc8341;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h230; din <= 32'hd7d46135;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02d; din <= 32'h7fa9b3e0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h321; din <= 32'hc4d3334d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h170; din <= 32'h258cccdd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d4; din <= 32'h7109253b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d3; din <= 32'h1ae53575;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ff; din <= 32'hcca6b2c4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14c; din <= 32'h09ea2867;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25c; din <= 32'h813f58a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h065; din <= 32'ha231db0c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h303; din <= 32'hf5c42dec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h123; din <= 32'h726784fe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h216; din <= 32'hca8c7b38;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08e; din <= 32'hca6c6c82;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35c; din <= 32'h0ea5b537;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h138; din <= 32'ha57e51e2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b8; din <= 32'hc3d08de1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h025; din <= 32'h3ee774da;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39b; din <= 32'hdb7255be;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h106; din <= 32'h4a4d5528;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h293; din <= 32'h94037dbd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h012; din <= 32'haceaf25d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h366; din <= 32'he8114167;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c1; din <= 32'hf6e74d59;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h239; din <= 32'ha9257db9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e6; din <= 32'h678e40c3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h335; din <= 32'h6cc0b362;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11e; din <= 32'h77aec888;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h203; din <= 32'hd625c641;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h068; din <= 32'h05348f52;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f5; din <= 32'h1581445e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13a; din <= 32'h6c685742;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d6; din <= 32'h816ef0bf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h011; din <= 32'h4af0fd4f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30d; din <= 32'h93edf082;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b7; din <= 32'h904db9da;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a5; din <= 32'he89acf52;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08e; din <= 32'h52d36f75;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h390; din <= 32'he1d276f3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d8; din <= 32'h54091070;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h231; din <= 32'h7875de35;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h026; din <= 32'hcdd529ac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h345; din <= 32'hb0c1883f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14f; din <= 32'h08553ec8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h262; din <= 32'h0491a22a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h019; din <= 32'habe33d1e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f0; din <= 32'hfad8e695;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14e; din <= 32'hfca2a846;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h258; din <= 32'he91fa34b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bf; din <= 32'h9c54a394;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3be; din <= 32'h2c04614b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h190; din <= 32'hf470a09f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h222; din <= 32'h8fd8fee0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0de; din <= 32'hcc818f44;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h325; din <= 32'hc5fea6ba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1eb; din <= 32'h89f2eecb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h223; din <= 32'h105b6484;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cf; din <= 32'hffdf9fd0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37b; din <= 32'h90cd0234;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h117; din <= 32'haf6be335;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cc; din <= 32'hb08ff40b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f0; din <= 32'h0d773dcb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h321; din <= 32'h7af6b374;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16d; din <= 32'he9129f6b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2dc; din <= 32'h2a56b33c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h027; din <= 32'hb16d35d5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fe; din <= 32'h973e077d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h145; din <= 32'h173a9ac0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26b; din <= 32'h7e4a21be;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h017; din <= 32'hadfaebcd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3df; din <= 32'h0c12231a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14c; din <= 32'h6fd205b3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cd; din <= 32'h33befab6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e1; din <= 32'h12fe29f8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fa; din <= 32'h57110390;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f1; din <= 32'h8ea854ee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h254; din <= 32'he4b28f15;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03a; din <= 32'h72f909df;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h351; din <= 32'h6143cacf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fb; din <= 32'h7a21cfcb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h246; din <= 32'h788e1b7c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ee; din <= 32'h9ae927dc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38c; din <= 32'h6602fa61;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h168; din <= 32'h002feece;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h269; din <= 32'h3a91451f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h059; din <= 32'h25ce3c6c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3df; din <= 32'he505d23f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h134; din <= 32'h52e7ed3a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26a; din <= 32'h5b495cf5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ab; din <= 32'h305ef27c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h358; din <= 32'hacd880b2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h179; din <= 32'h4f40d64e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f5; din <= 32'h6aa3492c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08f; din <= 32'hc535098b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f2; din <= 32'h404f8361;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ff; din <= 32'h396824a4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e7; din <= 32'hb86828eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0aa; din <= 32'h8f0169b0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h398; din <= 32'h0aaf4137;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h128; din <= 32'h0f9db5dd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e8; din <= 32'hf1209b92;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fd; din <= 32'hacc80d7e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h397; din <= 32'h24b26a0c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cc; din <= 32'h8915c68e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c2; din <= 32'h71989e82;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h053; din <= 32'h2ec8600d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h346; din <= 32'h0247a3b7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fb; din <= 32'h6862788e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h289; din <= 32'h4eeb0d1f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02a; din <= 32'hb8fffcbf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f2; din <= 32'h6dbb100f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cc; din <= 32'h78bc5ec6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e3; din <= 32'hb88d3844;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f3; din <= 32'hcf2a3b6a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38c; din <= 32'h124cbf84;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12c; din <= 32'h21e46a6f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h200; din <= 32'h261ba154;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fd; din <= 32'h13ea544f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30f; din <= 32'h0c40de04;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ef; din <= 32'hb4f06c04;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h297; din <= 32'h633f34f2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h065; din <= 32'h8e9d6b26;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35e; din <= 32'hc5812e73;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e4; din <= 32'hb1ef7bba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h290; din <= 32'h159c3863;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04d; din <= 32'he9811474;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33b; din <= 32'hd4de37fb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16e; din <= 32'h6a5bd5f2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28d; din <= 32'h0df6329a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h029; din <= 32'h6030d288;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h309; din <= 32'h0d0450ea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h164; din <= 32'hd330c793;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h214; din <= 32'hef80aea4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f0; din <= 32'hc007d37f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fd; din <= 32'h633a1b4f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c5; din <= 32'hb5408ee3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f1; din <= 32'h28666ba1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b6; din <= 32'h5afeea60;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h322; din <= 32'h3fe2db43;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h100; din <= 32'hd5822f80;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h220; din <= 32'hdde314e3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09a; din <= 32'h536f0cbb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h317; din <= 32'h460afb7e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18c; din <= 32'hab6d9dfc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h237; din <= 32'hb3e2c254;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h045; din <= 32'hb9195d43;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b0; din <= 32'had6f0204;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h158; din <= 32'h6dfe8e3d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f0; din <= 32'he1bb4c28;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ac; din <= 32'h6fb072ea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h336; din <= 32'h112f8491;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h121; din <= 32'h2e5f5594;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d1; din <= 32'heff1538e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0da; din <= 32'h696957ac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38f; din <= 32'h707ebbde;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c0; din <= 32'hf8ab33b8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h283; din <= 32'h42e17abc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h010; din <= 32'h96467dd2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h300; din <= 32'h332cd3c8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f3; din <= 32'hc18ec431;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h275; din <= 32'h9a263cd9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h007; din <= 32'h0f61409d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fe; din <= 32'h6b3f729a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h156; din <= 32'hd5088371;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29d; din <= 32'h03e75779;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09f; din <= 32'hf4f13c14;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fe; din <= 32'h849626a7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h137; din <= 32'hfc8d97d0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h287; din <= 32'h6797410d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03f; din <= 32'h3e3370a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3de; din <= 32'h87058a40;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h130; din <= 32'h62c52282;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h283; din <= 32'hed593c26;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fe; din <= 32'h690e5761;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d1; din <= 32'h0acd1950;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ee; din <= 32'h4dd8d89c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b0; din <= 32'hed584716;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h082; din <= 32'h306fec52;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h315; din <= 32'h1b4f6cd1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cf; din <= 32'h543c0392;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b4; din <= 32'h3513006e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h067; din <= 32'h30c1bd7a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h337; din <= 32'h63a0f35a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1be; din <= 32'hff3e6c74;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23b; din <= 32'h4c853203;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h001; din <= 32'hbc576a29;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3dd; din <= 32'ha6893ce4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h141; din <= 32'hbb0f1214;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c6; din <= 32'hdc26fb94;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h066; din <= 32'hde030baf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h343; din <= 32'h9b922cf5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12d; din <= 32'h45a0d871;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h296; din <= 32'hd9a4ceed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04f; din <= 32'h6c52482d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h348; din <= 32'h8a98806e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12e; din <= 32'hcac4863f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e7; din <= 32'h4d1685b8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h096; din <= 32'hc89a71fd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ff; din <= 32'hbb58fe99;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h174; din <= 32'he671cc0e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h236; din <= 32'h0e49297c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h059; din <= 32'h81ef0cca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h335; din <= 32'ha93baca9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12c; din <= 32'h1ccc28d6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d4; din <= 32'hdd04325f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f0; din <= 32'ha15c93a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38a; din <= 32'ha384af0b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h182; din <= 32'hc2b38f1b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28a; din <= 32'ha15f5b03;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02a; din <= 32'hc4614393;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h349; din <= 32'hb5d08e95;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h135; din <= 32'he6c1bb0c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f2; din <= 32'h0de8b796;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h017; din <= 32'hf599dc66;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ab; din <= 32'hd9a46823;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a5; din <= 32'h99ba31b4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2dc; din <= 32'hdf74dceb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h070; din <= 32'h4ecf4593;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39e; din <= 32'h1f7c3686;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h137; din <= 32'h3ed5cf1a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22c; din <= 32'h72fa5cd8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b9; din <= 32'h0e9239da;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31c; din <= 32'h38356947;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h120; din <= 32'h6c28bfb0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ab; din <= 32'h5f776bb2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04a; din <= 32'hf0f44b60;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35f; din <= 32'h57df8142;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e3; din <= 32'h2933eadd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ad; din <= 32'h751990c1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b3; din <= 32'h3db9aa18;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37c; din <= 32'h7af2de08;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b9; din <= 32'h52435322;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h206; din <= 32'hb29a0721;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h044; din <= 32'hf86d5f82;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34f; din <= 32'hc088ef00;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h183; din <= 32'h763e311e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a3; din <= 32'hdf6cf7de;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h045; din <= 32'h5062abce;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d9; din <= 32'hb7fb7950;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11e; din <= 32'hf7f8e532;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ca; din <= 32'h070939ee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03c; din <= 32'hf8c07677;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32d; din <= 32'h66ff1825;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h137; din <= 32'hfc8f41f6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c7; din <= 32'h3b1ee872;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h033; din <= 32'h13b37993;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c6; din <= 32'hff5b76be;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h100; din <= 32'hc79e1a5c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h261; din <= 32'hfadfc055;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c2; din <= 32'h7d09a6bb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e2; din <= 32'hafee5912;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c8; din <= 32'h08a2aec8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h257; din <= 32'hd52fd572;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h016; din <= 32'hd97a9a80;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bf; din <= 32'h3975e663;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c6; din <= 32'h38c3568d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h249; din <= 32'h14fe1021;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a1; din <= 32'hdbd085da;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h388; din <= 32'h5c7b9e45;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f3; din <= 32'h337082fa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d2; din <= 32'hb795cbd1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ed; din <= 32'h67eae2ba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cd; din <= 32'h345dbdec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h130; din <= 32'h5c67f9e2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h271; din <= 32'hbe681582;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f2; din <= 32'h8b90e661;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h308; din <= 32'h64ba7e7a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16a; din <= 32'ha6981d20;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h242; din <= 32'h4d6d2e23;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b2; din <= 32'hb33de6f3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f8; din <= 32'h2579c35b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16b; din <= 32'h3bdb6364;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h287; din <= 32'h48589055;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h020; din <= 32'h224ca55c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31a; din <= 32'h2ede3ce1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19a; din <= 32'h79d0a188;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h275; din <= 32'h8cdaa8d7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04c; din <= 32'hd5de3763;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d5; din <= 32'h204dcb4b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cc; din <= 32'h9de7f8d0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ce; din <= 32'hf90f8959;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e7; din <= 32'h7a2147b3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h397; din <= 32'h921eae78;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h127; din <= 32'he3e35ac0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28e; din <= 32'hcdea5487;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cc; din <= 32'hd4ab8cbf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h330; din <= 32'h47766fa0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15b; din <= 32'h9caeafe2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29d; din <= 32'h6ffa3bd6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07e; din <= 32'hf9923fc7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a0; din <= 32'h8efa25fc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h103; din <= 32'h30c70416;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h221; din <= 32'h3fff8633;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h085; din <= 32'h949674d3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38f; din <= 32'hc49410c3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c6; din <= 32'h7c83ccee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h287; din <= 32'hee641e85;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08d; din <= 32'hc18c2cf7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h332; din <= 32'hee72219a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h116; din <= 32'h8b7e3100;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29d; din <= 32'hb2542f6f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h014; din <= 32'hbb4e266d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38b; din <= 32'h35fdcba2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12c; din <= 32'h50225061;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25f; din <= 32'h76248361;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ba; din <= 32'hc432ff08;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h385; din <= 32'h6897f26a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ad; din <= 32'hde2a56b6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h200; din <= 32'hbc6b3619;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ce; din <= 32'heb457347;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h330; din <= 32'haad5f16a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16f; din <= 32'he55fcab2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2fb; din <= 32'h2ed32aba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ae; din <= 32'hd4b8d767;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h383; din <= 32'h167343e0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b9; din <= 32'h0de600f5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h234; din <= 32'h861665fd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f9; din <= 32'ha1713f94;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h300; din <= 32'h0e51f49c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ce; din <= 32'hf8d4c7a4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h233; din <= 32'h064cdc67;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03e; din <= 32'h0e928b7c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33c; din <= 32'h3f0abd48;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c8; din <= 32'hd47a0f42;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2cd; din <= 32'hab10fe51;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h068; din <= 32'h5d7d37f3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h361; din <= 32'h6abcd9b5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a3; din <= 32'h5e60bd0d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e9; din <= 32'h99b61bbb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e4; din <= 32'h48eb7894;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h367; din <= 32'h8b0b4cc7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bc; din <= 32'h5c1303b7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29c; din <= 32'h12e02c89;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e3; din <= 32'hfa25ad3a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h399; din <= 32'h62b06bfc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17e; din <= 32'hb485fdf7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22f; din <= 32'hdc3a133c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h077; din <= 32'h12d26b3d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h301; din <= 32'hb6e1fa40;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d1; din <= 32'h85c59b66;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f7; din <= 32'hcb55f6c5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07a; din <= 32'h3b77e732;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h372; din <= 32'h6684402d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h145; din <= 32'hea3cb8d0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a0; din <= 32'ha88d6741;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fd; din <= 32'h80faca98;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30e; din <= 32'h08f89a58;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15c; din <= 32'h81583c15;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h295; din <= 32'hdc7f19f3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bf; din <= 32'hc3a607d7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3db; din <= 32'hab52d3e6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h130; din <= 32'hc20ac350;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27a; din <= 32'h26178d85;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h091; din <= 32'hcc018340;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3da; din <= 32'habc905ae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ef; din <= 32'h25c8b499;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21c; din <= 32'h395a0130;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e9; din <= 32'hba7ee8b5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h314; din <= 32'h023279fe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ae; din <= 32'h039b98b2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c3; din <= 32'h7fad9394;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b3; din <= 32'hc4fa252b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34b; din <= 32'hd5796d17;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a4; din <= 32'h11c27f0d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e9; din <= 32'h94941587;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h070; din <= 32'h60602183;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h316; din <= 32'h5aed7da1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h110; din <= 32'hd0a9b884;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ba; din <= 32'ha98d8fd5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h014; din <= 32'h704a8592;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f8; din <= 32'hd6b0d68e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ec; din <= 32'ha6fc79c9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21d; din <= 32'hd79140ff;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h086; din <= 32'h3dd8a892;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h302; din <= 32'h5d4d9296;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a0; din <= 32'h8cd93379;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25b; din <= 32'hda1c2bd6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02e; din <= 32'h97da25ad;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h334; din <= 32'hfcdb65d1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h169; din <= 32'hc12f602f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24b; din <= 32'h670deec9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ca; din <= 32'h095da10b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32c; din <= 32'h93722e8f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h173; din <= 32'h0efe3719;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bd; din <= 32'hb75d1694;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h078; din <= 32'h30c44476;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h376; din <= 32'hdbb548a2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cc; din <= 32'ha9805d62;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h204; din <= 32'h7328376b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09e; din <= 32'h7be55711;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h320; din <= 32'h7cb86d34;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13e; din <= 32'h22234a6b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h204; din <= 32'h80e17e5d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h055; din <= 32'hfa7db9ac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a8; din <= 32'h96a460c0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h111; din <= 32'h126f4411;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e6; din <= 32'h3b7cb175;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00a; din <= 32'h094f7f95;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38a; din <= 32'h7298726d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15e; din <= 32'hb1cd33b6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d8; din <= 32'h56ac6efb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e2; din <= 32'h5aa10957;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3af; din <= 32'h32694b3c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h177; din <= 32'hbaf91e3b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b4; din <= 32'h037bcfec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e4; din <= 32'h0fe5df01;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d8; din <= 32'h22c23fce;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h105; din <= 32'hb9952040;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h261; din <= 32'had504bac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b7; din <= 32'h3431ad91;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30d; din <= 32'h44403255;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13a; din <= 32'h4c1cd2a5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28e; din <= 32'h78919d5b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04c; din <= 32'h868148e0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h335; din <= 32'h8132c674;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e7; din <= 32'h22bf7973;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29b; din <= 32'hafcf018a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05f; din <= 32'h36296ec6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3da; din <= 32'h5d77d963;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15b; din <= 32'hbf49e4c8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20a; din <= 32'he616bf3a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cd; din <= 32'h84babc62;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h391; din <= 32'hcb777e65;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17b; din <= 32'h63393a73;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h264; din <= 32'h07e2da43;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c2; din <= 32'hb72f7b89;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h317; din <= 32'h7f903e6c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h196; din <= 32'h4e18db9c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28e; din <= 32'hef097fbc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h031; din <= 32'ha15a6191;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32a; din <= 32'haffe2919;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h180; din <= 32'h4dbc4bec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c1; din <= 32'hcce00038;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h027; din <= 32'h583497fc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h380; din <= 32'hb274a29b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18e; din <= 32'hdcac3c83;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h208; din <= 32'h4818f799;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ea; din <= 32'hb64a1eaf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h300; din <= 32'h54387e4b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12d; din <= 32'h120cf93b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20b; din <= 32'h06ac418b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c0; din <= 32'h1daded4b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b5; din <= 32'h8a42fbc1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h107; din <= 32'hc251e4bf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23b; din <= 32'ha7b1a0af;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h010; din <= 32'hc58ebf29;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f4; din <= 32'h6ad63620;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h156; din <= 32'he45a820f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24b; din <= 32'h0c402c59;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h019; din <= 32'h222b9e1e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fc; din <= 32'h260e863f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h136; din <= 32'hcb8ffe0b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h239; din <= 32'h4ba23dd4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d7; din <= 32'h89468274;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a8; din <= 32'hf6c43437;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1dc; din <= 32'hc9dff92f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h266; din <= 32'he672614b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fa; din <= 32'h1d8079a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31c; din <= 32'h67467704;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15b; din <= 32'hd9529972;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a9; din <= 32'h083d2270;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0df; din <= 32'h157c570a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h346; din <= 32'h49cf885f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h133; din <= 32'hb877df68;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f8; din <= 32'hd25b8b77;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03b; din <= 32'h6546cbaa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bb; din <= 32'h0c0a2836;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13d; din <= 32'hc2f201d3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h216; din <= 32'h23ccd863;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h003; din <= 32'ha4048d4c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33b; din <= 32'h4b401855;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15b; din <= 32'h44eef548;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e3; din <= 32'h36102906;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ae; din <= 32'h740f93c6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3de; din <= 32'hbdfd5f8c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h158; din <= 32'h460fd770;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23b; din <= 32'h6cf1abee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h029; din <= 32'hffc7cbc8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h344; din <= 32'hc7b11f2b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14d; din <= 32'h13da26f5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h224; din <= 32'h710e4268;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h004; din <= 32'hca80ce5e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35f; din <= 32'h3be19e3a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h142; din <= 32'h5bea589e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22a; din <= 32'h8ca944ed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a5; din <= 32'hd8f4ccc6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h304; din <= 32'hfd2e0568;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h166; din <= 32'h12947123;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h234; din <= 32'h14bcd8c5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ea; din <= 32'h7d94ea50;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fd; din <= 32'h6828a372;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18d; din <= 32'h5cda8106;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e8; din <= 32'h079133a5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0af; din <= 32'hb59295d1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h396; din <= 32'h5ee1a9b4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h128; din <= 32'hbf034e6c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h274; din <= 32'h54b3a93a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h027; din <= 32'h3cfeb1d7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cb; din <= 32'h3f86aea7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14a; din <= 32'h3bf50240;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h214; din <= 32'h7414e9e2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h004; din <= 32'h0b0e445a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30f; din <= 32'h8ada87e8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h167; din <= 32'he720e085;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h253; din <= 32'h423c63eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f4; din <= 32'hfec460df;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h345; din <= 32'haf87c963;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h190; din <= 32'haee66104;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b0; din <= 32'hcb85bda8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ae; din <= 32'hdc7be8b6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h380; din <= 32'hcacae5c1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h182; din <= 32'h673da666;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h256; din <= 32'hb1e9737a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h017; din <= 32'ha5a8d7bb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35d; din <= 32'h2417710c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h148; din <= 32'h9aaaf61b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24c; din <= 32'h80c5e8fe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a3; din <= 32'hf83b3b94;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a9; din <= 32'h6851987b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18d; din <= 32'he1b0eb2d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h223; din <= 32'h503b5777;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h036; din <= 32'h5d174974;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39d; din <= 32'h646dc571;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h124; din <= 32'ha42d7180;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26c; din <= 32'hb47ef17d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h007; din <= 32'haa3fa564;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h308; din <= 32'h0b0895fb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d2; din <= 32'hf6db8871;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a4; din <= 32'h0d2f9336;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h048; din <= 32'h814f6952;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h394; din <= 32'h267e1d5f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16c; din <= 32'ha491692b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h260; din <= 32'h7b01821f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h026; din <= 32'h156e2ecd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cd; din <= 32'h76e2284a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16c; din <= 32'h2165de61;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a7; din <= 32'h266716f2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h051; din <= 32'h7de6e4ee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fa; din <= 32'he710f44f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h161; din <= 32'h2b7e9015;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h220; din <= 32'h1f4c41a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ce; din <= 32'hbe2679ba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ea; din <= 32'ha6899489;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h115; din <= 32'hbf5dd001;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h290; din <= 32'he46941e1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h039; din <= 32'hb3c205de;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35d; din <= 32'h3c566bc6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h187; din <= 32'h3c0624e3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h264; din <= 32'h4c2625c7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h097; din <= 32'h80247ef1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31c; din <= 32'h140210cd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18c; din <= 32'h97a695bd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e6; din <= 32'hc25cc8e6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h082; din <= 32'h9b185807;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h385; din <= 32'h098b1d93;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19e; din <= 32'h0dfd5d90;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e3; din <= 32'hd4967b94;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h019; din <= 32'h5a09d628;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h334; din <= 32'hda524f83;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h152; din <= 32'hda725e45;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2dd; din <= 32'h659371cb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h082; din <= 32'hee6e8ff9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ab; din <= 32'he6acfab5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12c; din <= 32'ha3fdf0e4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h247; din <= 32'ha75e6ee9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06d; din <= 32'h03d930e9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h306; din <= 32'h4dd563fd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h176; din <= 32'hec89d29a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h245; din <= 32'h7eee5fb3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f7; din <= 32'hb6fe2128;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h380; din <= 32'h11593c94;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19e; din <= 32'h687c7b5e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a5; din <= 32'h1ca95a40;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h030; din <= 32'h95bce7fc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b4; din <= 32'h1e65712d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a0; din <= 32'hd4d9773d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a3; din <= 32'hf4268779;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h042; din <= 32'h09bbaf9d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h324; din <= 32'hdca83893;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10a; din <= 32'h4b4ca048;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2dc; din <= 32'h20f32435;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h041; din <= 32'hc4326137;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35f; din <= 32'h5f5d3cc3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e8; din <= 32'h6f4bd0b8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h241; din <= 32'h2e746e2f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h032; din <= 32'hcc757eaa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h391; din <= 32'h038f1729;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h149; din <= 32'hf67179d5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24e; din <= 32'h52ecfdab;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h006; din <= 32'hc828aa95;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h333; din <= 32'haa0173f7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h132; din <= 32'hd55135bc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h264; din <= 32'ha1716aff;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h096; din <= 32'hdd9e6b44;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d6; din <= 32'h31eb0e13;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h199; din <= 32'he2afaa77;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29a; din <= 32'hf8660c1a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0bd; din <= 32'h10339599;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h306; din <= 32'h05953e23;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h146; din <= 32'h8584bad6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h23d; din <= 32'hffd4151f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a3; din <= 32'h3505fd76;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37a; din <= 32'h67beaf08;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14e; din <= 32'h00249eed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h272; din <= 32'h6a4a5ed2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e1; din <= 32'h59fd2ad2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32a; din <= 32'h246eaa62;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14f; din <= 32'h20640717;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h200; din <= 32'h6e3b8cd3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c6; din <= 32'h808e117e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b3; din <= 32'h0e3c1703;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h133; din <= 32'ha15fc5d8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h214; din <= 32'h694e87f5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09b; din <= 32'hff7aec36;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h373; din <= 32'h4c02cf07;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h179; din <= 32'hd57cc9e9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h276; din <= 32'h0e1f26bf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h092; din <= 32'hd960b561;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a6; din <= 32'h00f146c5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h182; din <= 32'h140bba5a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25b; din <= 32'h4c5fabcf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d0; din <= 32'h4d264c65;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e6; din <= 32'h93c1ef48;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19c; din <= 32'h2e1ef7a5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h270; din <= 32'ha8bbc216;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h038; din <= 32'h6859d373;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31e; din <= 32'h0c2a7b95;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h165; din <= 32'h2020bd2c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2dd; din <= 32'h87c16278;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fc; din <= 32'hb64bd24b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ae; din <= 32'he242c9eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f1; din <= 32'hb3a54ff0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29d; din <= 32'h4b5c1613;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h088; din <= 32'h5494e756;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a3; din <= 32'h21b8a186;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h121; din <= 32'h1f39897e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22f; din <= 32'h3c360bfe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a7; din <= 32'h285e720e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b8; din <= 32'h31b55bbf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19f; din <= 32'h6e3eb824;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h276; din <= 32'h8d9d4226;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08b; din <= 32'h1d0aebd1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h302; din <= 32'h90475fb5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d2; din <= 32'h1fee7044;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h228; din <= 32'hcd139432;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h077; din <= 32'hf2b73790;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h311; din <= 32'h12941d3c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cb; din <= 32'hf2a78cdd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h269; din <= 32'h7e448c90;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08b; din <= 32'hd074f239;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h386; din <= 32'h1bb213bb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1df; din <= 32'h566fed59;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d5; din <= 32'h42fcdcc3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07f; din <= 32'h6e1b8b43;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h301; din <= 32'h4f50386d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10b; din <= 32'hff3ece54;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h256; din <= 32'hba8fe543;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06d; din <= 32'ha6d27a62;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b3; din <= 32'h67bb7b0f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1aa; din <= 32'hbc8ecd55;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26a; din <= 32'h49e22018;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f8; din <= 32'h32561ecc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39c; din <= 32'h52081850;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h172; din <= 32'hf3852270;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h235; din <= 32'he0937b20;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04c; din <= 32'h92fd663e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d0; din <= 32'h17706dc1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h109; din <= 32'hbdf65c52;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h262; din <= 32'h9ea2d53b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a4; din <= 32'ha93389b3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b6; din <= 32'he94809d6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e1; din <= 32'hc50b9706;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28f; din <= 32'h83cb6415;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h094; din <= 32'h6b2f7a32;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37b; din <= 32'hfbd3568a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19c; din <= 32'h8867af9d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b6; din <= 32'h24e6dce4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09a; din <= 32'he95d2a8f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h331; din <= 32'hec4bef07;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c8; din <= 32'ha99a33b6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h292; din <= 32'he6cedb35;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d1; din <= 32'hc14f9ea9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a8; din <= 32'h2890c3f0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bf; din <= 32'h0242617f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21b; din <= 32'h01af28b2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h068; din <= 32'h3d02d73f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b7; din <= 32'h986f6703;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h152; din <= 32'h1e848b3f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f5; din <= 32'h44438416;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h002; din <= 32'h2c0d332e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h326; din <= 32'h8e434745;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10d; din <= 32'h1aef7c33;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bc; din <= 32'he1ad93e6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d3; din <= 32'h02c90187;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d0; din <= 32'h5dddacf7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17c; din <= 32'h9318c981;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h220; din <= 32'h41c081f4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h089; din <= 32'hc186befb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34c; din <= 32'h11a06eed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15d; din <= 32'h79a96449;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h275; din <= 32'h6aade938;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h014; din <= 32'h882faf63;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fa; din <= 32'ha093222a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fe; din <= 32'h07807f8b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h234; din <= 32'hf6cad3cf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f4; din <= 32'h85959c97;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d2; din <= 32'hde533ab9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1bc; din <= 32'h98a01fe2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h220; din <= 32'h279708c6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h065; din <= 32'h01d2def3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ba; din <= 32'h7a221fe0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h118; din <= 32'h61540dc0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h201; din <= 32'h97eb02da;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a4; din <= 32'h91dcc617;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h360; din <= 32'h3bf8a357;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f3; din <= 32'hcba4a836;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h262; din <= 32'hc4b3a1ef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h012; din <= 32'h755dd018;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h303; din <= 32'hcca72aee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h175; din <= 32'h9fe3e23c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f6; din <= 32'hf6a95fd5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02f; din <= 32'h1ffe8395;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d9; din <= 32'h82398903;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ad; din <= 32'hd9d98d08;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h293; din <= 32'h2ef5f3a4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h012; din <= 32'hdf6537bd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37f; din <= 32'hd48ac143;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h163; din <= 32'hc4777a9b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21a; din <= 32'had3330b4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h042; din <= 32'h33c730bd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38b; din <= 32'hb2b28df4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h144; din <= 32'hdef61138;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25d; din <= 32'h2328b7cd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h080; din <= 32'hb4a06f60;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38a; din <= 32'he9a39c25;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18d; din <= 32'hf552a542;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2da; din <= 32'hf15ceb3f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05b; din <= 32'h839f8818;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f1; din <= 32'h30600b93;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f4; din <= 32'h4bb8143d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e3; din <= 32'he02ff81a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h072; din <= 32'h2e799549;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h306; din <= 32'he620b889;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h115; din <= 32'ha9aa4a02;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f0; din <= 32'h4c73ddf2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h036; din <= 32'h36725405;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h336; din <= 32'hfcdafd8b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h170; din <= 32'hf645b48d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h29d; din <= 32'h90895cb2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h079; din <= 32'ha314fd4b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ba; din <= 32'hda98f207;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ea; din <= 32'h4596fa23;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d4; din <= 32'h0702d416;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h091; din <= 32'hc7613579;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h325; din <= 32'hd2f4ae86;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fa; din <= 32'h7f425bb1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h222; din <= 32'hde161ca1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fc; din <= 32'h41ecc37c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b2; din <= 32'h826c06a4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17c; din <= 32'h94f1a5bd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22f; din <= 32'h3cc786a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02f; din <= 32'hfdd2a710;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h336; din <= 32'hf1cf2171;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10d; din <= 32'h0c9de389;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a4; din <= 32'h811eba74;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f1; din <= 32'h2d8ae93f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a2; din <= 32'h27b53ce8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ff; din <= 32'hcc0e0115;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h281; din <= 32'h3677f7ec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h092; din <= 32'h4654ab20;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ed; din <= 32'h753faa97;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h153; din <= 32'h24eb2a9a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h224; din <= 32'h02f1a406;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h057; din <= 32'h468bd7c4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37a; din <= 32'hcf293110;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14d; din <= 32'h36d56bc8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h282; din <= 32'h1490dff7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06c; din <= 32'h9b716223;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h397; din <= 32'h6b6d833c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h134; din <= 32'h15dea278;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d9; din <= 32'hd3054d35;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09e; din <= 32'h6f5392c8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c2; din <= 32'hb1cb90e2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h145; din <= 32'hadc0cd6b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c4; din <= 32'h182b31ba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02a; din <= 32'h19c4bd18;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h340; din <= 32'h6627a32b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11d; din <= 32'h257007e7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c3; din <= 32'h7fefdb31;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h003; din <= 32'h5b0d72f6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ee; din <= 32'h1980416e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ce; din <= 32'h45764530;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bf; din <= 32'h5bd6b4cb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f7; din <= 32'h7d9d07b7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36f; din <= 32'h541522a4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h181; din <= 32'hda00f8d9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f1; din <= 32'h236a5d00;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h018; din <= 32'h375cc31f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h350; din <= 32'h25194c54;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h147; din <= 32'h55b6047e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h212; din <= 32'he826c285;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0af; din <= 32'h42565a4a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h354; din <= 32'h4760b74b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17b; din <= 32'he1b2523f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h244; din <= 32'h625e8f22;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h097; din <= 32'hd50d59df;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h364; din <= 32'h7e2fae97;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h121; din <= 32'hd5f28282;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d8; din <= 32'h8d4247ea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06a; din <= 32'ha60ae5b5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38b; din <= 32'h0655a4e5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h140; din <= 32'hb951ce02;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2db; din <= 32'h8782ec51;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ca; din <= 32'h3e331bb0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b1; din <= 32'h198111d2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18b; din <= 32'hce4a0bdd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f1; din <= 32'h189c6cfb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h008; din <= 32'hd9c53c5a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32d; din <= 32'h7ec7795c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h126; din <= 32'h6bf105e1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h203; din <= 32'hb47d55e7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b3; din <= 32'h981bfeaa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3da; din <= 32'h93b6dbaa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h152; din <= 32'h51d19833;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h247; din <= 32'h0340a5f6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h031; din <= 32'hbfb83dcc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h306; din <= 32'h833cfb08;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fc; din <= 32'h3ccc8899;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h272; din <= 32'h5252c4bd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04e; din <= 32'h0727dac3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39d; din <= 32'h9a594517;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11d; din <= 32'h383452a8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e3; din <= 32'he245c815;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cb; din <= 32'h0ff96ac9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h355; din <= 32'h6fe506e6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b8; din <= 32'hec04b8ed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20b; din <= 32'h57fb5e3c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06d; din <= 32'h59646204;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h314; din <= 32'h2fd830ef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ba; din <= 32'hcf612233;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2be; din <= 32'h916bd924;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h052; din <= 32'h4fc698df;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h396; din <= 32'hb800f33c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1c9; din <= 32'h9e88733f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21b; din <= 32'h90093977;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e8; din <= 32'h468de7a1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h331; din <= 32'h415a10f5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16a; din <= 32'hbdc3a880;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h227; din <= 32'h49a617b4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h008; din <= 32'h5358c663;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h377; din <= 32'hefeb48f0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h133; din <= 32'hdfb20e21;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26c; din <= 32'h1bd170f8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ef; din <= 32'h70df65f2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h339; din <= 32'h8d04855a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a4; din <= 32'h58d53b03;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f8; din <= 32'h38ffe23f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05f; din <= 32'h2f8b541c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h314; din <= 32'he9bcde8d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h102; din <= 32'h55634c64;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h220; din <= 32'h45d0e65d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h010; din <= 32'ha6f81d8f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h343; din <= 32'h9a0ccad0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h158; din <= 32'h6d272922;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h220; din <= 32'hbf7b72b8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h078; din <= 32'h32c9bcb0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30b; din <= 32'h17a600ae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1db; din <= 32'h58bf9b5e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d9; din <= 32'h2b3aa22d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0da; din <= 32'h951402de;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h305; din <= 32'h77c5fdc1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13d; din <= 32'h4662067a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b0; din <= 32'hb1d4f5e1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c8; din <= 32'h592e2cd9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h380; din <= 32'ha826dcfb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11d; din <= 32'h706bfa11;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2df; din <= 32'h33f8f941;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h058; din <= 32'h39498d4b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h337; din <= 32'h795e057c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1fd; din <= 32'h20bcf404;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ef; din <= 32'h33514cb8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c8; din <= 32'hb1e6a3a9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h326; din <= 32'h7f64097e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16e; din <= 32'hfc496298;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2fc; din <= 32'h52d80e64;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b5; din <= 32'h9232db84;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h320; din <= 32'hafd919ad;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h12a; din <= 32'ha3c8342d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h266; din <= 32'ha121d7a0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h035; din <= 32'h88003c9d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ac; din <= 32'h36aa2ea1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b1; din <= 32'hdeed2606;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b8; din <= 32'h9bdd099d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b5; din <= 32'hfbd90163;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f8; din <= 32'ha7ec6303;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1aa; din <= 32'hc815af78;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28b; din <= 32'h55e25369;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03e; din <= 32'h57d5ab20;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e9; din <= 32'h6bab3271;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h152; din <= 32'hc5f3a1cb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c3; din <= 32'h69f115a7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h095; din <= 32'h4fed08d2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3dd; din <= 32'ha503d739;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h170; din <= 32'h0eb3e1e3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20a; din <= 32'h2fb43951;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0aa; din <= 32'haa769199;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38d; din <= 32'hc22eea05;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h137; din <= 32'h2f53c538;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f6; din <= 32'h2b5d7115;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h020; din <= 32'h72aa1123;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h361; din <= 32'h704806e1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a1; din <= 32'h9a4bd4a1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b1; din <= 32'h8f0ab588;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06a; din <= 32'h61667edc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h334; din <= 32'h99e53ff6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1be; din <= 32'hf45e0457;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h255; din <= 32'haf8296ac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h006; din <= 32'ha3f9314d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h339; din <= 32'h865ae23d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h165; din <= 32'h9845d0ea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h239; din <= 32'h1f057b5d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0aa; din <= 32'h2bf2c2c6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h360; din <= 32'h7f61967d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13b; din <= 32'h3ea5842d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27b; din <= 32'hbdb0bac3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f9; din <= 32'h64751ff2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h390; din <= 32'hd69b421e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e7; din <= 32'hca4629bf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2da; din <= 32'h63d0d021;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h083; din <= 32'h398f437c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38d; din <= 32'h28841fed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1ad; din <= 32'h90a8849a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h248; din <= 32'haae826e6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h017; din <= 32'hbc228a4c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33e; din <= 32'hea4a5c11;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h131; din <= 32'h416ebf52;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bb; din <= 32'hdfa76244;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d7; din <= 32'hb7c13ac1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bc; din <= 32'h370cdf54;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h13b; din <= 32'h0cb5799f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h256; din <= 32'h02f15dd9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h019; din <= 32'he4f21cd5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ac; din <= 32'h5aee3df0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h136; din <= 32'h43d838d5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24d; din <= 32'ha86901cf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05a; din <= 32'h0379c9a8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a8; din <= 32'h10ddf66d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17a; din <= 32'h9df374bd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h266; din <= 32'h5dc2fc32;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f0; din <= 32'h27a2c2ca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33f; din <= 32'h5c7a5e4f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h15b; din <= 32'h4508e94f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22c; din <= 32'h59f91ac0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h067; din <= 32'hdf5a8fd9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31f; din <= 32'h1cb1f79d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h196; din <= 32'h33a33e8c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ce; din <= 32'h6f23b07b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0df; din <= 32'ha00a8784;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ac; din <= 32'h13b0f780;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h188; din <= 32'h0194c005;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h253; din <= 32'hb1ec9a41;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07b; din <= 32'h5b3f8440;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37b; din <= 32'h30984f43;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1e3; din <= 32'he1c744e1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20a; din <= 32'hd0422d31;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0df; din <= 32'hb6df7452;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h371; din <= 32'h9416ce82;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cc; din <= 32'h8c6f8e6f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h263; din <= 32'h8740dec0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ef; din <= 32'hde5d2320;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ab; din <= 32'h0c639b5c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14c; din <= 32'hc7b11f90;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d5; din <= 32'hfbe9ccf6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h074; din <= 32'h40e69305;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3cb; din <= 32'hf7704529;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d8; din <= 32'h393c44f7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h250; din <= 32'he28d105f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cb; din <= 32'he1565e8a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d2; din <= 32'heaccf2b9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h160; din <= 32'hed68c729;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h20b; din <= 32'hac9979a9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h039; din <= 32'h698af5f6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39c; din <= 32'h99c324f8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f5; din <= 32'h69e6af08;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a2; din <= 32'hcafbf8aa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h083; din <= 32'h2a39d807;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37d; din <= 32'h2d79accc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h153; din <= 32'h1c5497df;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a3; din <= 32'hb226724a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h010; din <= 32'h0c893a51;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b0; din <= 32'hbfc29871;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h157; din <= 32'h892cd3ec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2be; din <= 32'hf10821fa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h089; din <= 32'h64a54327;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h349; din <= 32'h8209a9b8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18f; din <= 32'h72d746e8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h256; din <= 32'h47b87b91;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c0; din <= 32'ha9e70d13;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38d; din <= 32'h849dedc5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h10a; din <= 32'h12820a7d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d5; din <= 32'h040af2a5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04d; din <= 32'h837a0dec;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h362; din <= 32'h74f2907e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cb; din <= 32'h491518c3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h212; din <= 32'h904801c5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h089; din <= 32'hffb86f57;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f5; din <= 32'h22be9b13;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h191; din <= 32'h064991cc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e1; din <= 32'heeb7c347;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09a; din <= 32'h1ae3e9ca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c8; din <= 32'h914da0df;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h165; din <= 32'habc03986;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e9; din <= 32'h04ba6361;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h051; din <= 32'hac31eeb5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a4; din <= 32'h1420daaf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1eb; din <= 32'h6f935fc1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e6; din <= 32'h7d3fab48;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01c; din <= 32'hb0ed73e1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h396; din <= 32'h4cbaac90;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h187; din <= 32'h5303fd7b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22c; din <= 32'hda637656;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h021; din <= 32'h91a841ac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h346; din <= 32'h5104f77b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19e; din <= 32'h1ee34de4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a1; din <= 32'h647c8021;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h027; din <= 32'he6a6cd84;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30f; din <= 32'h3e549ea7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17f; din <= 32'h38a9e93d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2ce; din <= 32'h6a8d1c4f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h076; din <= 32'h77487bc8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h374; din <= 32'hb278604d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h182; din <= 32'h3e27a7e8;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h21a; din <= 32'h7c7368b2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04a; din <= 32'h03b4060b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39a; din <= 32'ha3d35987;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b6; din <= 32'h9dd174c7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h278; din <= 32'hefd9aebe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h044; din <= 32'h4993f44a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33f; din <= 32'hd7092189;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h19f; din <= 32'ha54ba5f3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h239; din <= 32'ha117d9a7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0fa; din <= 32'hecd60f69;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34d; din <= 32'h8bb9ed43;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h123; din <= 32'hfc241392;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h247; din <= 32'h3338debe;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h029; din <= 32'h9edc88c2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h388; din <= 32'hba05cae9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16a; din <= 32'h900e2877;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h254; din <= 32'h419ba710;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h095; din <= 32'h29457092;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h338; din <= 32'h32506796;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16d; din <= 32'h4232b214;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h238; din <= 32'hcd7cfb45;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09e; din <= 32'h8e52c5e9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c8; din <= 32'h1ac0a083;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h178; din <= 32'hac2dcd5f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h233; din <= 32'hb53d0fa7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cd; din <= 32'ha82f5707;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b1; din <= 32'hb62982db;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h174; din <= 32'h815a9881;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2b6; din <= 32'h9a9baa3c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f6; din <= 32'h00bcd8ae;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h320; din <= 32'h9144e463;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h17f; din <= 32'h8491a6eb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h215; din <= 32'h2a580011;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e1; din <= 32'h1921ee26;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h388; din <= 32'hc8e30f82;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h151; din <= 32'h36ac7d20;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c6; din <= 32'he394b877;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h056; din <= 32'h9ad78601;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c7; din <= 32'h2cc9402c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b8; din <= 32'h95c7b25a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2bd; din <= 32'h462572e2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h060; din <= 32'h06f19059;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ab; din <= 32'h70fefaf6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h148; din <= 32'h051584dd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h222; din <= 32'h6a2d3dfc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0ac; din <= 32'h0ae7cd36;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h384; din <= 32'ha978cfce;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h107; din <= 32'h121a919a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a1; din <= 32'h3541917c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f8; din <= 32'hf0cea937;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h368; din <= 32'h703fed34;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h133; din <= 32'h8d9661aa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25a; din <= 32'hbb940572;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e1; din <= 32'hc423b472;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bb; din <= 32'ha8cd7687;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h122; din <= 32'hc1bc9374;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h216; din <= 32'he7edfa13;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cb; din <= 32'h52912d30;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d3; din <= 32'h4a2c5553;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h180; din <= 32'h5feecf59;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27f; din <= 32'h7121a655;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b7; din <= 32'h4223025d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39a; din <= 32'h0127e358;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16d; din <= 32'h7d971c4d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h217; din <= 32'h8844500c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02f; din <= 32'h9328af6b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ff; din <= 32'h8895e4b4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f8; din <= 32'h6d3c8da3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2fd; din <= 32'h1df6c73b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05a; din <= 32'hd4d5e665;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h392; din <= 32'ha6beaa65;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h16b; din <= 32'h1eb2a11c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h27e; din <= 32'he5e931bd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h02c; din <= 32'hf547fd91;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36d; din <= 32'h6d3c198c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h112; din <= 32'h91bbd148;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h218; din <= 32'hf1298beb;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01e; din <= 32'h69f3f9ee;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38b; din <= 32'h21516de5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1d6; din <= 32'hfa83834d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h214; din <= 32'h901f3741;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h04f; din <= 32'h567cee84;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a4; din <= 32'hcd5dc748;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h130; din <= 32'h4c37a3ac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24d; din <= 32'hbc622ded;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06c; din <= 32'hdda92d2f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b5; din <= 32'h51c5f2a4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h123; din <= 32'h9cc4363f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h226; din <= 32'ha035a5c1;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0df; din <= 32'h4096c56d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h337; din <= 32'h8b0947cc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h165; din <= 32'h37ddcf22;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d9; din <= 32'h8e4d0a36;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c0; din <= 32'h135b4a2d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a3; din <= 32'h539df8da;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1dc; din <= 32'h5ca2ae1d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c1; din <= 32'ha149d828;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h034; din <= 32'h843b2c2c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3fc; din <= 32'h4790dc34;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1b3; din <= 32'ha7e67a88;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h24a; din <= 32'h2b1c14aa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h061; din <= 32'h69b46a63;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34c; din <= 32'he22e902f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h185; din <= 32'h1f9ab84c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h250; din <= 32'he8a090e3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a5; din <= 32'hefd0aa92;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d2; din <= 32'h157d26ef;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18a; din <= 32'h12f3b95e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a0; din <= 32'h84e80c72;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b2; din <= 32'h611a193c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h328; din <= 32'h56f84998;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h121; din <= 32'h186aa143;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25c; din <= 32'h96110c3c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cb; din <= 32'h0606e201;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h347; din <= 32'ha56ce176;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h106; din <= 32'h0db1ec17;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h298; din <= 32'ha39a2bb3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00f; din <= 32'h1b7bae53;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h33b; din <= 32'h28120765;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h119; din <= 32'h75da3312;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h210; din <= 32'hfbc04c25;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h058; din <= 32'h9049553f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h32a; din <= 32'h14ebdea6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h194; din <= 32'h9d76f1a4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f5; din <= 32'h2fae2d42;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h046; din <= 32'haf72f47a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h332; din <= 32'h72d1c8d4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1f4; din <= 32'ha90e6877;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h273; din <= 32'h76f9681a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03a; din <= 32'h0739a9ba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3a5; din <= 32'h6774c4ac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h195; din <= 32'hce428c19;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h253; din <= 32'h16ee3f01;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00a; din <= 32'h12485460;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38a; din <= 32'h51cb66a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h169; din <= 32'hc1bae1e3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e2; din <= 32'hf8f89c0d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e9; din <= 32'h61b3e674;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3dd; din <= 32'h4d631029;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18e; din <= 32'h320c1845;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h28f; din <= 32'h951abbe5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00a; din <= 32'h0e47b8a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h366; din <= 32'ha17ae3b5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h18f; din <= 32'h712a0660;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c1; din <= 32'hdacbb633;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09b; din <= 32'hdd692816;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h356; din <= 32'hc07baf83;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h196; din <= 32'h431a4f6c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f8; din <= 32'h9656cc28;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h072; din <= 32'h4b2507d3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h386; din <= 32'h1da42748;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h120; din <= 32'h6c635a75;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h237; din <= 32'hc3d54171;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05e; din <= 32'hd492de44;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3dd; din <= 32'h960f6d04;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h197; din <= 32'h701e7240;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2e7; din <= 32'h5b7d1861;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e0; din <= 32'h62999a78;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ab; din <= 32'hcb384932;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cc; din <= 32'hfae07548;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h224; din <= 32'h3bc8a97e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01e; din <= 32'hb5e8f12d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h38d; din <= 32'ha636f31f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h11a; din <= 32'h5475db84;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2d8; din <= 32'h51ff67c9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d9; din <= 32'hc7b2edd9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37a; din <= 32'he87cab01;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h189; din <= 32'h1b47e3c6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h22e; din <= 32'h3c0a5465;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h069; din <= 32'h9db26d06;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e7; din <= 32'hcf76d29d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h108; din <= 32'ha7fa4f87;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h26f; din <= 32'h7dc387d9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h061; din <= 32'hbd22173b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bd; din <= 32'h1edfadbc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1cf; din <= 32'h80ff75b4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2db; din <= 32'hc6e41269;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00d; din <= 32'h898f9c90;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h381; din <= 32'h82490325;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h1a5; din <= 32'h726ecd02;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f6; din <= 32'hb2dca2ed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h043; din <= 32'h4fa8d5c3;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h382; din <= 32'h46d8ef90;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h150; din <= 32'hebaec8f0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2a8; din <= 32'h55e1d6a6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h09d; din <= 32'h9493aecd;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b7; din <= 32'h2496c498;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h174; din <= 32'h3b2e9bb9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h210; din <= 32'h3730921f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c2; din <= 32'h2b035201;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h368; din <= 32'h37964e18;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h14f; din <= 32'h7ebc2763;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2c8; din <= 32'h13a0c693;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h071; din <= 32'h4052e5ad;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h323; din <= 32'h2485b69b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h251; din <= 32'hc06a76c9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h052; din <= 32'h8e132fa5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bb; din <= 32'hf6b2709e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h292; din <= 32'h771dd79e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03f; din <= 32'h4cf42de2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h330; din <= 32'h009c5013;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h25c; din <= 32'h68015e14;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00a; din <= 32'hb9d35663;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31c; din <= 32'hc24df40b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h2f1; din <= 32'h318e11ea;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a8; din <= 32'h1137d06f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c7; din <= 32'hfec891c5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h299; din <= 32'hb6870590;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h043; din <= 32'h8f5fd326;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bf; din <= 32'h3f3d4d7e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h292; din <= 32'h3559825f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0c8; din <= 32'habd4844d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h313; din <= 32'h2f3be430;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b1; din <= 32'h6d88140f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3dc; din <= 32'h54c0a5d2;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07e; din <= 32'h0ef6f417;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c1; din <= 32'hc24b88de;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0e4; din <= 32'hd79c9bdc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h390; din <= 32'h39559784;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h01d; din <= 32'h4dff408c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h39e; din <= 32'h7e960249;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a2; din <= 32'h4c340f64;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3e9; din <= 32'hf39b2012;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f4; din <= 32'h740f305c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h312; din <= 32'ha16423a5;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h072; din <= 32'h0022d7b0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h324; din <= 32'h49df6447;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b2; din <= 32'h7ff4ad92;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3f2; din <= 32'h7447c69f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0db; din <= 32'h9750b7dc;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ba; din <= 32'h93d3bd05;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h05a; din <= 32'h94b23fd7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h317; din <= 32'h7903683b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h004; din <= 32'h1bd9c89a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h336; din <= 32'hf673fd1a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h037; din <= 32'h93ac6f94;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h37f; din <= 32'h14c91cde;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h08f; din <= 32'h0439b6c6;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h369; din <= 32'h366ee48a;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h082; din <= 32'hf0178b58;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h31c; din <= 32'h298e38bf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h089; din <= 32'h586cc080;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h388; din <= 32'hb8b8c5c4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h00f; din <= 32'h16566da0;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h30d; din <= 32'h2f69a973;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h092; din <= 32'hcedbef22;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3ae; din <= 32'hce62d958;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h03c; din <= 32'h1508c34e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h383; din <= 32'h7e23aae4;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h016; din <= 32'h8e92e5ca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h351; din <= 32'hc1934335;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0dc; din <= 32'h300b3aba;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h344; din <= 32'h83f68886;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d1; din <= 32'h964dacc9;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h369; din <= 32'hb7ef6c9e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h06d; din <= 32'h47abf80d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h302; din <= 32'hc1fece69;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0d2; din <= 32'h38f2f259;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h34a; din <= 32'hb0810a48;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h084; din <= 32'h47b5fb48;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b3; din <= 32'h349ce52c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h095; din <= 32'h8404fc88;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d2; din <= 32'h1a4e964e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07c; din <= 32'h332edb20;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h332; din <= 32'h4e1c80ed;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0a9; din <= 32'h3ef67f0f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h300; din <= 32'ha137a35c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f2; din <= 32'h2a179a53;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h35a; din <= 32'hca7e4340;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h007; din <= 32'h373b9fcf;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h347; din <= 32'h365835f7;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0f2; din <= 32'hc303db1c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3b0; din <= 32'h091aadca;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h054; din <= 32'hde35257d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c1; din <= 32'h3b453867;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h024; din <= 32'h5fc1350d;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3bc; din <= 32'hd1b0265b;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h099; din <= 32'h9de21880;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h302; din <= 32'h4e579068;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0b2; din <= 32'h0b2e49ac;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h338; din <= 32'h1ed41b8e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h074; din <= 32'h8ba27207;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h398; din <= 32'hc1605f77;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h036; din <= 32'hf5e32e67;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h342; din <= 32'h7cd0e83f;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h003; din <= 32'h8c3bb645;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3d5; din <= 32'h3ec7108c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h068; din <= 32'hb5c22f56;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h393; din <= 32'h091ba266;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h075; din <= 32'hd2eb190e;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h36a; din <= 32'h755392aa;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h0cf; din <= 32'he5d60368;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h3c1; din <= 32'hb894ca7c;
        @(posedge clk); en <= 1; wen <= 1; addr <= 10'h07a; din <= 32'h1eb54d25;

        // Finish
        @(posedge clk); en <= 0;  addr <= 10'hxxx; din <= 32'hxxxxxxxx;
        repeat (5) @(posedge clk);
        $finish();
    end

    always #1 clk = ~clk;
endmodule
