`timescale 1ns / 1ps

`ifndef INSTR_MACROS
`define INSTR_MACROS 1

`define NO_INSTR 2'b00
`define WRITE_INSTR 2'b01
`define READ_INSTR 2'b10
`define MOVE_INSTR 2'b11
`endif

module testbench #(parameter DATA_WIDTH = 32, parameter BYTE_ADDR_WIDTH = 8, parameter BANKS_ADDR_WIDTH = 2);
    reg clk;
    reg rst;
    reg [1:0] op;
    reg [BYTE_ADDR_WIDTH+BANKS_ADDR_WIDTH-1:0] addr;
    reg [DATA_WIDTH-1:0] din;
    wire [DATA_WIDTH-1:0] dout;

    inspec uut (
        .clk(clk),
        .rst(rst),
        .op(op),
        .addr(addr),
        .din(din),
        .dout(dout)
    );

    initial begin
        $dumpfile("waveform.vcd");
        // $dumpvars(0, testbench.uut.rst, testbench.uut.op, testbench.uut.addr, testbench.uut.din, testbench.uut.dout);
        $dumpvars(0, uut);

        // Initialize
        clk = 0;
        rst = 1;
        op = `NO_INSTR;
        @(posedge clk); rst <= 0;
        @(posedge clk);

        // Autogenerated code        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d4; din <= 32'h2ea53750;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h079; din <= 32'hed401f46;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h36e; din <= 32'h677a618f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h323; din <= 32'h97725dda;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3dd; din <= 32'h5b6a354c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a4; din <= 32'h4d318ca7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h385; din <= 32'hf17b0f5c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h15f; din <= 32'hefa460e5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h011; din <= 32'h3b81d309;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ad; din <= 32'h61d1a67f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h25c; din <= 32'he110fb4e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h36e; din <= 32'hdcfc5948;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22f; din <= 32'h08fc791d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h163; din <= 32'he75eab93;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h158; din <= 32'h4b6a5db0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h34d; din <= 32'h8fa1552c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2dd; din <= 32'h40480720;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c0; din <= 32'h6a07536b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h154; din <= 32'h75a3e386;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ed; din <= 32'hca791052;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h249; din <= 32'hcd11921a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h11a; din <= 32'hb9925d22;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h110; din <= 32'h3600c35a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2cc; din <= 32'h1395eefe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h125; din <= 32'he33afe96;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d9; din <= 32'hd39176ec;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h03b; din <= 32'h09851351;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h363; din <= 32'hede893c4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h13c; din <= 32'h25298b93;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b2; din <= 32'h29260d69;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ca; din <= 32'hc88b25cb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h205; din <= 32'hb75d1114;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d8; din <= 32'hc9650928;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h146; din <= 32'hf14d6230;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h197; din <= 32'h880120c2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f9; din <= 32'hac629ed6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f8; din <= 32'hdac90f34;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1cf; din <= 32'h7360eb24;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3eb; din <= 32'hf6900bb2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ca; din <= 32'h7eb120fb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h335; din <= 32'hd5c1d6f4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e9; din <= 32'hb1cdc3e4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d4; din <= 32'h8462371d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b2; din <= 32'h731f5840;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h11a; din <= 32'h7d3d8966;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f9; din <= 32'h72ac2c00;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b9; din <= 32'h2fe61b7a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3aa; din <= 32'h8a7c70b8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16b; din <= 32'h81190019;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h225; din <= 32'he9f8d9c2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h245; din <= 32'h7df01ea4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h224; din <= 32'hc038e65b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h317; din <= 32'hc880412b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h27c; din <= 32'h40d7de8e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f5; din <= 32'h797d4d2c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h004; din <= 32'h6c15d3c3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2eb; din <= 32'h6c740849;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h208; din <= 32'hde229936;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e0; din <= 32'hb20e54d0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d8; din <= 32'had75f58a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h28b; din <= 32'h71db22e6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a1; din <= 32'hdd65fe17;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h366; din <= 32'h852ca88a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ce; din <= 32'h451b5351;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h29d; din <= 32'h9ccd3903;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h159; din <= 32'h6a5314df;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h232; din <= 32'hb2eeb293;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d4; din <= 32'hc5e7f978;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h167; din <= 32'h55914099;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1bf; din <= 32'h6924e99f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h29a; din <= 32'hd6eec1cd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h17b; din <= 32'h13cf53dd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16b; din <= 32'h45ceec21;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h176; din <= 32'hcd240b7a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h28a; din <= 32'h9209c009;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h12a; din <= 32'hc7da917d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e1; din <= 32'h66dd260f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f9; din <= 32'ha61abc97;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e4; din <= 32'hac863e19;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h208; din <= 32'ha9f221a9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h27e; din <= 32'hde7eecda;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1fd; din <= 32'h8bfc3045;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d3; din <= 32'h6c00a387;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1cc; din <= 32'hd05bdaed;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h384; din <= 32'h02cc2f70;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d9; din <= 32'h852af0bb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38a; din <= 32'h6d82dc0b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h19c; din <= 32'hec5c0aba;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h153; din <= 32'h47fcb4f8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d1; din <= 32'hc5011099;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00d; din <= 32'hc723ba28;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h373; din <= 32'h4d8a804d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e0; din <= 32'h4ae70b60;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h28e; din <= 32'h6d02a4d1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h107; din <= 32'h87317958;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a8; din <= 32'h0098d7c7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d3; din <= 32'h0ab5a06a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08e; din <= 32'h8d0d7d60;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18a; din <= 32'habd8b399;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h313; din <= 32'h3308c29a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b6; din <= 32'hb78f5b68;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h03c; din <= 32'h5191d242;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e0; din <= 32'h3d74fe74;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h325; din <= 32'heae0db6b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h080; din <= 32'hb123e2a6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b0; din <= 32'h81581390;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ba; din <= 32'h4a973fea;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h118; din <= 32'h6e6438da;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h33e; din <= 32'hd3490d3b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h029; din <= 32'h306f0767;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c5; din <= 32'hc72dbcda;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h09a; din <= 32'h2ef6440a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ed; din <= 32'h72c2701d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23b; din <= 32'h32d2f981;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h310; din <= 32'h52437e9c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h363; din <= 32'h36a1c9b5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h201; din <= 32'hb0d25b67;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37a; din <= 32'hcec4d824;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h290; din <= 32'h492aa2da;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h04e; din <= 32'he9fc339b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e4; din <= 32'h660ba8ba;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h017; din <= 32'hb8584830;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h229; din <= 32'hc0f0906b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h192; din <= 32'h2d381954;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ff; din <= 32'h1ee91e65;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h287; din <= 32'hb6cf8d52;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h29e; din <= 32'h70168c83;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h123; din <= 32'hb2c32a5f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h29c; din <= 32'h79798c38;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h012; din <= 32'h0a8a1b39;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1cb; din <= 32'h2e43528d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h251; din <= 32'h4f7e9029;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a7; din <= 32'hc587afed;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h264; din <= 32'hc0f181be;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h238; din <= 32'h341fd0a1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h143; din <= 32'hc8cd4815;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a8; din <= 32'hd028c5e2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ce; din <= 32'h879aace4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h299; din <= 32'hc0eb4827;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h282; din <= 32'h2ba74def;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b8; din <= 32'h6dff5d71;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h001; din <= 32'hb4192ea5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2aa; din <= 32'hc12b49fc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h359; din <= 32'hbc1b72e5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f7; din <= 32'hf926efbb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h27a; din <= 32'h6d0b3165;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f8; din <= 32'h972deb0e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h375; din <= 32'h959e591d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38e; din <= 32'ha59933df;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h26d; din <= 32'hb78e1113;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h343; din <= 32'hfd2582f9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h32d; din <= 32'h5a7402ba;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h261; din <= 32'h728a6c77;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h186; din <= 32'h3a002224;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08e; din <= 32'he98e9d0e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31c; din <= 32'h54439ef3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b3; din <= 32'he59cf326;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c1; din <= 32'hd5a5e9ca;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23a; din <= 32'h0fd4d89c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f8; din <= 32'h21405c1a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h316; din <= 32'he7245a0b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f9; din <= 32'hd548b064;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h065; din <= 32'h9986ff4e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3af; din <= 32'ha2778b9e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ba; din <= 32'hd62caa5e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h343; din <= 32'h6848977d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h191; din <= 32'h9d85440b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f2; din <= 32'hbb791c7a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2fe; din <= 32'h976fda67;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h12a; din <= 32'h4b1a022f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h038; din <= 32'hd637d58a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h06c; din <= 32'h1ae06344;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b1; din <= 32'h4a30962a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d1; din <= 32'h1287a62c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h297; din <= 32'h684ed1fa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ae; din <= 32'hf3d032e6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h317; din <= 32'heac0aad9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h390; din <= 32'h39f6feae;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h28a; din <= 32'hab05d620;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37c; din <= 32'h37f605ff;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h107; din <= 32'h15ced2cb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h26d; din <= 32'h5c1212ae;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38c; din <= 32'hc8727b00;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3eb; din <= 32'h1b48d141;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h125; din <= 32'h940716b9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h200; din <= 32'h1d8a23b8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ee; din <= 32'h94485c36;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f5; din <= 32'h106432bf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2bf; din <= 32'ha0cd5a58;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2aa; din <= 32'hbdd17f13;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h270; din <= 32'h5b56ec60;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0bd; din <= 32'h51a52012;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f9; din <= 32'h755a26b5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b7; din <= 32'hf9351829;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ce; din <= 32'hd30595a7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h20c; din <= 32'he40da49c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0de; din <= 32'h29360697;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h32b; din <= 32'ha6e40d7e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h016; din <= 32'hec18e2bb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e6; din <= 32'h8718c03b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h356; din <= 32'h5f943449;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h130; din <= 32'hf69d2675;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h335; din <= 32'hc3958529;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e4; din <= 32'h0bb4ec4d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b8; din <= 32'h381eb6de;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h041; din <= 32'ha1e9e3cb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h314; din <= 32'h4ae48acb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h075; din <= 32'h69953356;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h342; din <= 32'h0811f40a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h368; din <= 32'hcf0d4869;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1af; din <= 32'hf10c83c3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ea; din <= 32'hd62cc66f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h271; din <= 32'h837daa37;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1db; din <= 32'h7c030564;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b8; din <= 32'hac9a684c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h350; din <= 32'h27b15365;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h164; din <= 32'h312d104e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h035; din <= 32'hc58e40a2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h25d; din <= 32'h348436a4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c6; din <= 32'hdd501fca;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h157; din <= 32'h00908f5e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e2; din <= 32'hd54b212a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h350; din <= 32'h9eda545a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h189; din <= 32'ha0e30900;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31e; din <= 32'h9b6c82be;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h156; din <= 32'h8c7a1071;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f3; din <= 32'hd1fa3e35;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h370; din <= 32'heb194240;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31c; din <= 32'h2f8f4e9d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h225; din <= 32'h39b7be3f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08b; din <= 32'hc23cf73e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e5; din <= 32'hc48d0fbd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h36c; din <= 32'h0a9ad7ff;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h320; din <= 32'h5aed4ebf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38e; din <= 32'h7e738276;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d4; din <= 32'hbf7b30af;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08f; din <= 32'h402ff613;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ab; din <= 32'h9b4040ef;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h04b; din <= 32'h4b9de373;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h068; din <= 32'hc6972591;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e0; din <= 32'h7b04350c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h004; din <= 32'hf80b2e3a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h333; din <= 32'he426848d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2fe; din <= 32'h310e8456;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31d; din <= 32'h6df1c28f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f3; din <= 32'h43bbe7f7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c9; din <= 32'h2f6781b4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h30e; din <= 32'h6266b386;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h050; din <= 32'hc5828ca8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h008; din <= 32'h65167ea8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h24e; din <= 32'hbb3dcb9f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22c; din <= 32'hff27a71e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h044; din <= 32'h41957ac4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c6; din <= 32'hb3685aa6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f4; din <= 32'ha9382b5f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h372; din <= 32'h7daba396;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c1; din <= 32'he484de2f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f5; din <= 32'hb8cbc7eb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h171; din <= 32'hc21bcf2e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h257; din <= 32'h28d031d7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h068; din <= 32'h987052b7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2fb; din <= 32'h28bb56f9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h19d; din <= 32'hf054597b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h32c; din <= 32'h2a318943;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d9; din <= 32'he2975a10;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h311; din <= 32'h13cef648;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h34c; din <= 32'h6319d8e6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h053; din <= 32'h5cf1bee0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h344; din <= 32'he4b073d0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h223; din <= 32'h0ec6d260;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h06a; din <= 32'h519f15b0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h031; din <= 32'h04db436e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b2; din <= 32'hc93c9b02;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h24d; din <= 32'hf93e4677;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b2; din <= 32'he026c9be;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h211; din <= 32'h4bd6a9f0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h129; din <= 32'h9419e890;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h02b; din <= 32'h6ffec0fe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1fd; din <= 32'hb88fc589;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38b; din <= 32'hb5b18131;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h037; din <= 32'hc8e54e4d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h34d; din <= 32'h5609addb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h088; din <= 32'h67245517;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f9; din <= 32'hfc9d9741;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h244; din <= 32'h06e693f0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h020; din <= 32'hd536f0db;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h396; din <= 32'h4c6708b1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h11c; din <= 32'h5609c85c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h013; din <= 32'h2c5e12b5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16a; din <= 32'h06db46df;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ba; din <= 32'h489a503f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h268; din <= 32'hecc38a12;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h074; din <= 32'h5946f7e9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h03f; din <= 32'hd87c5cf1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h041; din <= 32'h899abb43;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e6; din <= 32'hc3a85328;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h355; din <= 32'he604163d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e4; din <= 32'h57715371;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h03d; din <= 32'h01c2648b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h07b; din <= 32'h0470f5bc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ca; din <= 32'h663393b3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h350; din <= 32'h28993a04;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h27d; din <= 32'hae3e5f2f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h371; din <= 32'h0d9b54b8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h380; din <= 32'h7b70d4eb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e1; din <= 32'h2fa8c24a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16a; din <= 32'h161384ff;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h157; din <= 32'h04b275d3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ac; din <= 32'h9cb46fe0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h30d; din <= 32'ha1e5aee9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23f; din <= 32'h610c9821;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18b; din <= 32'h23051229;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c2; din <= 32'hd52d6f26;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c4; din <= 32'h8a72bca0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h26a; din <= 32'h600ad7bd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3eb; din <= 32'hed5d46c9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f2; din <= 32'h31b252a1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h373; din <= 32'hc3f0c505;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h336; din <= 32'h5733948d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h24d; din <= 32'h916632ec;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h228; din <= 32'hef5e9aad;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h27d; din <= 32'h6351b88a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h175; din <= 32'haa20b0a3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h09c; din <= 32'hcdd64527;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h09f; din <= 32'hf5fc8e42;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h24d; din <= 32'h2c9e245d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h13c; din <= 32'h7406df9d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2cd; din <= 32'h3f0009f8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h270; din <= 32'h46f7d753;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h28d; din <= 32'h7e69f70a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h070; din <= 32'hd09f5c92;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0db; din <= 32'hdb8b4027;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h257; din <= 32'h959160a4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h061; din <= 32'h02e415da;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1db; din <= 32'hda6ab8e3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h160; din <= 32'h8c719514;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h315; din <= 32'haf5177b8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2a2; din <= 32'h93070107;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c2; din <= 32'hd165a0fd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h008; din <= 32'h36e0db52;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b2; din <= 32'h054c6a4d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h316; din <= 32'h552c1d5c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h197; din <= 32'h20b68fbe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h178; din <= 32'h3746ca86;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h290; din <= 32'h18af35d7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h29a; din <= 32'h0860b2db;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e3; din <= 32'h99029200;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1da; din <= 32'hb07e4bec;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h288; din <= 32'h196c627f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h310; din <= 32'hf37e23bf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h210; din <= 32'hd6502701;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a4; din <= 32'h01f0824d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h180; din <= 32'ha6fcd139;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h079; din <= 32'h9228f648;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h285; din <= 32'hf217843b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h372; din <= 32'h8d2aeed9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h028; din <= 32'h6e80cae7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h189; din <= 32'hcd369af2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0cf; din <= 32'h422baad4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h329; din <= 32'he0113ea3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h115; din <= 32'h7f3ed4d4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h186; din <= 32'hf3588679;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c2; din <= 32'hd168d541;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h297; din <= 32'h56045d10;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h26d; din <= 32'h747b18c9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2cd; din <= 32'h84c9a1b3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h124; din <= 32'ha7b9b5c2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2a6; din <= 32'hfb543f90;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h25a; din <= 32'hfe4cbe87;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ac; din <= 32'ha1167e6c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38f; din <= 32'h1a59f4d1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08a; din <= 32'h8e7fa93f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d7; din <= 32'h2fad8d09;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h057; din <= 32'h8ecf2d3c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a4; din <= 32'hda151f23;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h11f; din <= 32'ha00938b3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1af; din <= 32'h62eeb4a2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h19e; din <= 32'h23761e94;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22d; din <= 32'h41660a01;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h06a; din <= 32'h418e28a1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ac; din <= 32'ha011fce4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3dc; din <= 32'hca1a250a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d8; din <= 32'he98017b5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h368; din <= 32'hd5482c32;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h02c; din <= 32'h85f049ea;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h013; din <= 32'hf6109899;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h342; din <= 32'h9527b529;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b5; din <= 32'hb6a3c32b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1dd; din <= 32'h5de5cf82;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23e; din <= 32'h45a84ab7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18d; din <= 32'he3138e68;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3bc; din <= 32'h1001a536;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h25b; din <= 32'hb9b0135a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h188; din <= 32'h48792e68;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h072; din <= 32'hb9e000ba;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31c; din <= 32'hb01c5077;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h026; din <= 32'h9f3c93dc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h345; din <= 32'hd6d05d37;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h110; din <= 32'hf6d93573;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e5; din <= 32'h9302dc39;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h263; din <= 32'ha8aebd09;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h07a; din <= 32'h3fbdfd3e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16f; din <= 32'h539f1d11;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h069; din <= 32'h0b9cea7d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e2; din <= 32'hc0e37185;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h185; din <= 32'h25f065a9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e1; din <= 32'ha7beb252;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h054; din <= 32'ha8ed12da;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a9; din <= 32'h5c8ff059;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h168; din <= 32'h3850a25d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h11f; din <= 32'h2219b264;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d3; din <= 32'hf8d319d6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h04a; din <= 32'h943e5a8c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h05e; din <= 32'h4d0c1b87;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h188; din <= 32'he20bbf10;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ec; din <= 32'h836f8878;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ff; din <= 32'h90ddb5de;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h080; din <= 32'h3f43a996;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h170; din <= 32'h2f24b1a6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16a; din <= 32'hff9b463b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ea; din <= 32'h09687ff1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h177; din <= 32'hf637d5f2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h20c; din <= 32'h595a229e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d0; din <= 32'h5edbca2c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h240; din <= 32'h85b795b6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h20c; din <= 32'ha91c3926;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h145; din <= 32'h9dce6165;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1bf; din <= 32'he4dca4eb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h365; din <= 32'he071b094;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h159; din <= 32'h7ba2dbcd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h21b; din <= 32'hefc4cf62;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h12a; din <= 32'hcae4e590;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d0; din <= 32'hca5a10b4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h183; din <= 32'h7a02e9e7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h359; din <= 32'hcc590071;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h067; din <= 32'h1ce15a65;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h32e; din <= 32'h8b10973a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e2; din <= 32'he1d96747;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a4; din <= 32'hffb7b81a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h223; din <= 32'h5f636520;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23e; din <= 32'h3c383c28;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h088; din <= 32'h94f9363a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h276; din <= 32'h423bcd90;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f7; din <= 32'hb3a5cfe2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e8; din <= 32'h3e67e14c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2cb; din <= 32'hf161587a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e2; din <= 32'h594538c8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h371; din <= 32'h79572104;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b2; din <= 32'hefac28c3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h272; din <= 32'h0e96dc37;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c0; din <= 32'h3208e145;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d6; din <= 32'h434576a8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h059; din <= 32'h0de94f49;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3eb; din <= 32'h4fa86e38;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h095; din <= 32'h729b8b00;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h076; din <= 32'haa60baac;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h108; din <= 32'h68526fa5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h302; din <= 32'ha05ef898;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e4; din <= 32'hd205f494;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h27c; din <= 32'h6f67cd14;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h248; din <= 32'h7cdd8dfa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ac; din <= 32'h2c32b50a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ef; din <= 32'heaf22d80;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h35d; din <= 32'h1cb22add;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h145; din <= 32'h135766b2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1aa; din <= 32'hfa9b0213;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0bd; din <= 32'hc6d75b0d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h19a; din <= 32'hcfc98327;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f4; din <= 32'ha76325ca;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f5; din <= 32'hc3566398;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h27e; din <= 32'haa3f8bd8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h228; din <= 32'h7ca0bfaa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h20c; din <= 32'h8f043b82;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c4; din <= 32'h36a4e221;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b7; din <= 32'hb064bd1f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0db; din <= 32'h984fb135;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h048; din <= 32'hda3e76b5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h036; din <= 32'h9d6395a9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h09b; din <= 32'ha7bcec12;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h349; din <= 32'h6a4305ca;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h305; din <= 32'hb77efaa6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h06b; din <= 32'h01e187af;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h382; din <= 32'h62289ac9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h012; din <= 32'he9f67bbb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e4; din <= 32'h9a315e75;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b0; din <= 32'h2c3dded2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f0; din <= 32'hd2653f0d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h14e; din <= 32'h0cb91401;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h357; din <= 32'h2a4f19a3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h002; din <= 32'h3e276a16;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h160; din <= 32'h78a1326d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f3; din <= 32'h3da5cd42;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h203; din <= 32'hd5c7344f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2cb; din <= 32'he817be2c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22d; din <= 32'h26fc19b9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h046; din <= 32'h6b90ff3f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h297; din <= 32'hefdde4f1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h110; din <= 32'h70f2164b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c2; din <= 32'h3bcd8d12;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d7; din <= 32'h494f4bea;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h11b; din <= 32'hd6f350c7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h19f; din <= 32'hccdaab25;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e7; din <= 32'hd4643b2e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0fe; din <= 32'h861fae1d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b1; din <= 32'hc3dd96aa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h279; din <= 32'hdacf6348;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22c; din <= 32'h0382e3f6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h242; din <= 32'hbecd2539;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h392; din <= 32'h44249aa5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h350; din <= 32'h4906cd05;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ed; din <= 32'hdbdb0e3a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2dc; din <= 32'he8fec568;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h17a; din <= 32'hefcf12a2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22b; din <= 32'h5d06077f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2fc; din <= 32'hda5323a4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h015; din <= 32'h681be124;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f0; din <= 32'hd8cdeb13;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a3; din <= 32'h0bba4f4b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h213; din <= 32'h8bae8ab2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h257; din <= 32'h2e7471cf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h237; din <= 32'h69c87fde;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h128; din <= 32'h44eb4b4b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2dc; din <= 32'h3adfc53c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h077; din <= 32'h9821207a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1dd; din <= 32'h8ae962c0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ba; din <= 32'h699577f3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f5; din <= 32'hd5b0c898;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h364; din <= 32'h81aad768;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f2; din <= 32'h1ace7958;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3cd; din <= 32'hb8fe0d8d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00c; din <= 32'he99fc92a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h033; din <= 32'hcf72fe61;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ba; din <= 32'h7fe7e6d8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37c; din <= 32'h6ca14844;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ca; din <= 32'hb4a4ec2d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h30d; din <= 32'h23ea9509;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h15a; din <= 32'h20e5ebd3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2be; din <= 32'h4ffc993a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h252; din <= 32'h2248b5f9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h062; din <= 32'h66351a8d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h091; din <= 32'h8ef694b6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h307; din <= 32'h97aac21b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ab; din <= 32'h6ad3826c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h388; din <= 32'haa7fa66c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h27e; din <= 32'hc55fbac3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b3; din <= 32'hd2c2c2b8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ef; din <= 32'h8b379b7f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b0; din <= 32'hff81c425;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h169; din <= 32'h4756b4ae;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b3; din <= 32'h2a6bb866;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2eb; din <= 32'h3dddd0bd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h335; din <= 32'h1ffa9fff;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1de; din <= 32'h0491ee7c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h050; din <= 32'h5b6d8389;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f1; din <= 32'h0e99d6cc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h26d; din <= 32'ha16f39dc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h357; din <= 32'h38119054;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h074; din <= 32'h26914457;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d6; din <= 32'hbad6a122;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b8; din <= 32'h4f59300a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h36d; din <= 32'h388a0f0e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h148; din <= 32'h185f4f2b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h06c; din <= 32'hc9a568da;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ad; din <= 32'hf3637970;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h027; din <= 32'h09230ab6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h072; din <= 32'h1eb22cca;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38e; din <= 32'hea132ce3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h342; din <= 32'hf141d77d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h05d; din <= 32'h0dc20e4f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h11c; din <= 32'h641b2324;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h32e; din <= 32'h366365f5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h33c; din <= 32'h60c6f3fb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h052; din <= 32'h158c2548;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h21f; din <= 32'h9103de8a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h354; din <= 32'h92014fce;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h337; din <= 32'h34967b22;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h255; din <= 32'h5b952baa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38f; din <= 32'h9709212c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f7; din <= 32'h85ce29c3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2cd; din <= 32'hae6fd117;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h207; din <= 32'h0b9ca345;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h089; din <= 32'hbe5c3058;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e6; din <= 32'h08533cfe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h089; din <= 32'h9bb5db4a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h05a; din <= 32'h02a8bc86;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c2; din <= 32'h69651ef6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ae; din <= 32'hd629550b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h191; din <= 32'h7686a0cc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h253; din <= 32'hd13e54e4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c8; din <= 32'heac9d4a4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e1; din <= 32'h7a80b2a7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3db; din <= 32'h843e1973;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f8; din <= 32'h0f9c8b89;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h214; din <= 32'h752ccb97;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c7; din <= 32'hc1f2c0e9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e0; din <= 32'h9c806008;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b3; din <= 32'h46465f91;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d9; din <= 32'h9dd14742;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h191; din <= 32'heb283ae7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h380; din <= 32'h291be88e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b6; din <= 32'h4031d41a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h116; din <= 32'h088ec7aa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h041; din <= 32'h8b373be0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h155; din <= 32'haec06687;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h254; din <= 32'he8f75183;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h32d; din <= 32'h3e9b2254;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h305; din <= 32'h2900feba;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h312; din <= 32'h1bc19980;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h116; din <= 32'hcc426653;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31d; din <= 32'hfbd7b97d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f1; din <= 32'hc2202f88;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h024; din <= 32'h7c7087db;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h132; din <= 32'hf80cc3e3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h203; din <= 32'h3ac64941;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08f; din <= 32'h1668045f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e0; din <= 32'h2208dcc0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h193; din <= 32'h8048553f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ff; din <= 32'h33635c3f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h350; din <= 32'h34e8061e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h212; din <= 32'hda468710;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ba; din <= 32'hfb2242ee;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h196; din <= 32'hfe53fdce;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e3; din <= 32'h2c31ecb9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e2; din <= 32'h3eb405c0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22b; din <= 32'h2ba2629b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a1; din <= 32'h022d69bb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h307; din <= 32'h9ec2bcbc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a3; din <= 32'h65ea31ab;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b8; din <= 32'h65edcb69;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08a; din <= 32'h75b98797;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h098; din <= 32'h724da128;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ba; din <= 32'h673eb895;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d4; din <= 32'h51461a06;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2a4; din <= 32'ha75c6816;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h109; din <= 32'he85a6480;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1de; din <= 32'hbea03eb6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h354; din <= 32'h555ead22;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h213; din <= 32'h0157c60b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h26b; din <= 32'h17dc3a4c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h033; din <= 32'h64f895a5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h397; din <= 32'h8e9977b2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h349; din <= 32'hf9280a81;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a9; din <= 32'h22f6a7fb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ee; din <= 32'hf0870f54;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00a; din <= 32'h09ce85bb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h098; din <= 32'habf5ce56;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2fd; din <= 32'h6f72a2fd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h291; din <= 32'had3ec2c1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1bd; din <= 32'h757fee1f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1df; din <= 32'h09500fc9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h025; din <= 32'h48cf1cd0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c0; din <= 32'h42da82ef;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h329; din <= 32'h92ed341e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3bc; din <= 32'he3f57bfd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h06c; din <= 32'h70179004;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h196; din <= 32'h0108f9de;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2a1; din <= 32'h74f79fde;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a9; din <= 32'hefed0597;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a0; din <= 32'h9be3193b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c1; din <= 32'h600d0545;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h02d; din <= 32'h3993ec02;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b8; din <= 32'h7f85f831;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h097; din <= 32'h0c271df1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b2; din <= 32'h8dbaf279;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h087; din <= 32'h6cd6f28f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h366; din <= 32'h1968eb45;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b3; din <= 32'h81712337;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h20c; din <= 32'he142d95a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c7; din <= 32'h922fb543;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h039; din <= 32'h8b5b3945;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h089; din <= 32'hff581fe7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ac; din <= 32'hcacb1826;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ae; din <= 32'h99983340;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h067; din <= 32'h6894078e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22e; din <= 32'h358c2f6b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e0; din <= 32'hc9906e98;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0df; din <= 32'hde9818d4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c6; din <= 32'h9922538e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c7; din <= 32'hf5348bc8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a2; din <= 32'h10ead638;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08d; din <= 32'h148e93dd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f1; din <= 32'h30994a22;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2a1; din <= 32'hcf90b166;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h376; din <= 32'he95b52cd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h242; din <= 32'h228a4677;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3cf; din <= 32'h1c20844c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h28a; din <= 32'hef1349ec;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f1; din <= 32'h6d64faa3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ba; din <= 32'h28a4860e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h07b; din <= 32'hae281857;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h26f; din <= 32'h1c75f104;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h328; din <= 32'h016848e3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h21a; din <= 32'h66388a3d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h372; din <= 32'he167470d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h289; din <= 32'h894cbadd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h21f; din <= 32'hc2c74818;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h216; din <= 32'h3484bc96;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h158; din <= 32'hcc2812c8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h047; din <= 32'h7c7100d8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h173; din <= 32'hb5c382d0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1fb; din <= 32'he7673db5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h078; din <= 32'h1bdca3d5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h09a; din <= 32'h19868bcf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h20f; din <= 32'h09cf3456;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ea; din <= 32'h17fc6a17;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d8; din <= 32'hc46236a1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h058; din <= 32'haab6a8fe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e0; din <= 32'h2a2f881f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h091; din <= 32'h39b75d13;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d1; din <= 32'h5836e304;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h004; din <= 32'h75d20778;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f3; din <= 32'habb415bd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h017; din <= 32'hc3a45f58;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h268; din <= 32'h93f192df;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h303; din <= 32'h3c28c6db;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1dd; din <= 32'h85b73f6b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b8; din <= 32'h5ffee634;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37a; din <= 32'ha5772666;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h286; din <= 32'h5fc75c0b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h116; din <= 32'h6dd38b80;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ee; din <= 32'h459a9129;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h216; din <= 32'hbee6506f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h298; din <= 32'hfd057de1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3fd; din <= 32'h4d0ad7d9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h306; din <= 32'h1b77a040;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h069; din <= 32'h25cea02b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b2; din <= 32'hdeb27bdd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f9; din <= 32'h66f206c0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h361; din <= 32'h047957d1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h216; din <= 32'hc65c4e71;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h097; din <= 32'hfe1a68ce;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h058; din <= 32'h61191b70;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h163; din <= 32'h8ca599aa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h294; din <= 32'h66419095;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a5; din <= 32'hb289fd7d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c0; din <= 32'h81e18667;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22b; din <= 32'hc53fc5a2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b2; din <= 32'hd9bcec7f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h04f; din <= 32'hc14d6c2e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c8; din <= 32'h6052d8b9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d3; din <= 32'hebb4f742;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h393; din <= 32'h8576c72a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h03f; din <= 32'he1c92c27;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e3; din <= 32'hab41a6f2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h375; din <= 32'h0dc6a738;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h24d; din <= 32'h42adfd22;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h016; din <= 32'h42e93df7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h35a; din <= 32'h7dd9a1fe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h15a; din <= 32'ha4e6f517;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h159; din <= 32'h6a8d9a6e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h35e; din <= 32'h17c9096c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h186; din <= 32'h70ed04c3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h124; din <= 32'h6f55b79f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38f; din <= 32'h0c5a9bea;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16b; din <= 32'h87d4b4a4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h20a; din <= 32'h9afd07e6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e4; din <= 32'h24b38439;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ef; din <= 32'h9df683e4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h220; din <= 32'h16d3580e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d2; din <= 32'ha549bd2c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h21e; din <= 32'hbc7aac82;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h296; din <= 32'h19e2c60a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h390; din <= 32'h846656b2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c9; din <= 32'h1421d7fb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h10c; din <= 32'hc31e9ae6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h39d; din <= 32'h483658a2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h107; din <= 32'he5acb8c3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h169; din <= 32'h8a0d018c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h074; din <= 32'h62bf6021;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3dc; din <= 32'h7419bf2a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h03f; din <= 32'hfc71993d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h12c; din <= 32'hbeb8a22f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e2; din <= 32'h3cb63a56;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22d; din <= 32'he0d8c9fa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c1; din <= 32'hc869cdf7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h165; din <= 32'h8af80a96;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h275; din <= 32'hbf0feb87;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f1; din <= 32'h15460470;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h25d; din <= 32'h254642d2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h105; din <= 32'hf6f18b33;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e7; din <= 32'hb4a006bd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c5; din <= 32'hb6479f48;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h159; din <= 32'hac1247de;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2a1; din <= 32'h9a39ccfb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h35f; din <= 32'hf9f05757;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c9; din <= 32'h908c06cd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a0; din <= 32'hd210da5a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h313; din <= 32'hff6ca76a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b8; din <= 32'h7d2d183c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b2; din <= 32'hc5a4170a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b0; din <= 32'h08fcd929;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ef; din <= 32'h3fd78dd2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18c; din <= 32'h552f1680;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37b; din <= 32'hcc132575;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18e; din <= 32'hab916372;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h308; din <= 32'h9ecef5e0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h115; din <= 32'hc4baa5b9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h05f; din <= 32'hbeefbfba;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ea; din <= 32'hdba13705;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2fc; din <= 32'ha9aae899;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3fb; din <= 32'h27ef3a44;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d7; din <= 32'hbe7c1304;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h318; din <= 32'h82995f9c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c9; din <= 32'h16bd4b6c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e9; din <= 32'h10179ff8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e0; din <= 32'haa0242d9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h165; din <= 32'hff995482;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e1; din <= 32'hdea79cc8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a1; din <= 32'hd889b0cb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h25f; din <= 32'h852334cf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h12a; din <= 32'h1a293941;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2fb; din <= 32'he35b5b2f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e9; din <= 32'h1b271763;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h024; din <= 32'hb39cd23d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37b; din <= 32'h39657217;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e3; din <= 32'h4ac31c4a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b3; din <= 32'hcc3cb987;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c8; din <= 32'h7de66463;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18f; din <= 32'h43bf4e11;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h036; din <= 32'h1e210fa2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h309; din <= 32'h30958c83;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1fd; din <= 32'h81e0059b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d1; din <= 32'h4e40c612;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h324; din <= 32'h73e88005;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37d; din <= 32'h1b0c81f9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ee; din <= 32'hc6ccc45e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ad; din <= 32'h3c24000e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h04d; din <= 32'h612535c2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h36b; din <= 32'h2ae90a1d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h196; din <= 32'h07bb2466;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h045; din <= 32'h2bc866e5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h345; din <= 32'hea409f48;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e8; din <= 32'h018a6deb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1cf; din <= 32'hcb80697c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h11e; din <= 32'h512becfb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h028; din <= 32'hecca6205;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2be; din <= 32'h3b4188da;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e1; din <= 32'h2962d771;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h152; din <= 32'h0e3c3cc7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h02f; din <= 32'hd813cf52;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h010; din <= 32'hee1a5466;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h180; din <= 32'h5fc34a0a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h393; din <= 32'ha5a709a1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f1; din <= 32'he7ea9bb8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h181; din <= 32'hf2ccaf4b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c3; din <= 32'h4597ab12;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h14b; din <= 32'hd422baa4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0de; din <= 32'h8710be10;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ad; din <= 32'ha2375530;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h300; din <= 32'h5fac5332;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e2; din <= 32'he5282f4f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h382; din <= 32'h6c09e522;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h33c; din <= 32'h4c4bdc00;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d5; din <= 32'h46b6127e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h349; din <= 32'hc5291a02;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h27c; din <= 32'h899dc771;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0aa; din <= 32'h062da442;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h236; din <= 32'hcd779745;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h042; din <= 32'hc7b86b9c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h295; din <= 32'h7230aef0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h347; din <= 32'hb0518652;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b8; din <= 32'h07e87d8b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h235; din <= 32'hce393917;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h06f; din <= 32'hd2638c04;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h04c; din <= 32'h3613715f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h07b; din <= 32'ha5858e8f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h35b; din <= 32'h6b0c8928;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0bd; din <= 32'hf6043f30;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f0; din <= 32'ha7a5c520;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b0; din <= 32'h1a7f53d4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h236; din <= 32'h651c7155;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0fd; din <= 32'h97c83c35;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h32e; din <= 32'h6179beea;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h076; din <= 32'h84959cc7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e7; din <= 32'h96e56213;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h099; din <= 32'hcb345126;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h278; din <= 32'h1992a722;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e7; din <= 32'h650b9e1c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0bb; din <= 32'h7d02e807;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3df; din <= 32'h2c3e517e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f5; din <= 32'hd5fde961;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h004; din <= 32'hc04f61f5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h04b; din <= 32'hc8f616ee;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22d; din <= 32'hfa313581;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h117; din <= 32'hf30edc83;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ba; din <= 32'he618439b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2bf; din <= 32'h7c83c59e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b5; din <= 32'hd995a6eb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h206; din <= 32'h9945fdff;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e2; din <= 32'h00868659;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h055; din <= 32'hd50548cb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b8; din <= 32'h60bc009c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h03a; din <= 32'h69f16aca;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h054; din <= 32'hfb42fd84;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00d; din <= 32'ha4b19206;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h022; din <= 32'hfc9befa4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h13f; din <= 32'h35e189b1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h155; din <= 32'h858eeae2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2fb; din <= 32'ha339c20e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1da; din <= 32'haa023864;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h053; din <= 32'hefcb4416;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h39d; din <= 32'hc396a80a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h168; din <= 32'h6763a0aa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e6; din <= 32'h4aed5c1e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3fe; din <= 32'h6a570498;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h193; din <= 32'h0ffe0ad5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18c; din <= 32'h6fe37481;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h256; din <= 32'h6bbdde15;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h113; din <= 32'h04069fa2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1da; din <= 32'hdd2e7ea4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h068; din <= 32'hc66b7c33;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h329; din <= 32'h5deff75e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h341; din <= 32'h0feb1ac0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c7; din <= 32'hfd798690;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3df; din <= 32'h32c29fae;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h26a; din <= 32'h79031137;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h327; din <= 32'h3bdbd8b8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h012; din <= 32'he0a9c963;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h146; din <= 32'ha353c36c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h359; din <= 32'hc225327a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3dd; din <= 32'h866fc350;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h337; din <= 32'h3722f5e5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f8; din <= 32'h79dd8381;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h281; din <= 32'h832cca4d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h134; din <= 32'h597592d8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1fb; din <= 32'h9574c93d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h003; din <= 32'h85c87224;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f5; din <= 32'hf43a9fe1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d0; din <= 32'he9cd700d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h394; din <= 32'hf083cd99;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h107; din <= 32'h6da0ff11;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h389; din <= 32'h61e3a04b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c4; din <= 32'h01c7719d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e7; din <= 32'h675a7e29;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h092; din <= 32'hf01ea36e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h159; din <= 32'h48935c85;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1cf; din <= 32'h35554475;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h023; din <= 32'h2ae5dbe3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22a; din <= 32'hdb97f88e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3fe; din <= 32'h3a7fcf90;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3da; din <= 32'h0bc53a43;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h187; din <= 32'h4dbb531a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h135; din <= 32'h47560316;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h331; din <= 32'hc7f698cd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1fd; din <= 32'h3a3cab0b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h07c; din <= 32'hb094ffac;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h164; din <= 32'he17bf220;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c7; din <= 32'h23016ea5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h194; din <= 32'haf641d80;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h030; din <= 32'hdbdb2473;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h258; din <= 32'h96fce18c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d1; din <= 32'ha7d92e37;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b7; din <= 32'hc4d618ac;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1dd; din <= 32'ha05b5497;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h055; din <= 32'hd652098c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3cf; din <= 32'h93280d9c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00b; din <= 32'h2da2feef;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0db; din <= 32'hbbe75532;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e0; din <= 32'hfd1d89ea;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h277; din <= 32'h72d8efea;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h256; din <= 32'h9aa4cbd0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h35d; din <= 32'h5af23a55;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h168; din <= 32'h1321e0fa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h02b; din <= 32'h1683727b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h052; din <= 32'hb6f7868b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h12b; din <= 32'h23534114;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f8; din <= 32'hca191fe4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18b; din <= 32'hd32b715a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h181; din <= 32'h12cff594;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h365; din <= 32'he26341e0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h36d; din <= 32'hb7fce032;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37d; din <= 32'h2acea6f3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08b; din <= 32'ha4045081;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b6; din <= 32'h5e0829f7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d5; din <= 32'h0b648d97;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2cf; din <= 32'h8c6c17f4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h01d; din <= 32'h9058598f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b7; din <= 32'h2622a533;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h212; din <= 32'h1b534438;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h057; din <= 32'h4e5ba382;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h17a; din <= 32'he986a394;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b9; din <= 32'h2d88a075;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b2; din <= 32'h08f1ebb9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h305; din <= 32'hc072262e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h065; din <= 32'hccddfd7d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h279; din <= 32'he553f7f0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h10f; din <= 32'hcde86944;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h04d; din <= 32'h594ecd59;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h063; din <= 32'h7cc3c1d7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3db; din <= 32'h19d929b0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f1; din <= 32'hf159ead4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3fa; din <= 32'hbea47bf0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h321; din <= 32'hec3b365d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ad; din <= 32'h2f50df02;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h259; din <= 32'h09bc7fec;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h39c; din <= 32'hf80f096b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f0; din <= 32'h5f29401b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h264; din <= 32'h46777c23;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h020; din <= 32'h92b7b254;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h24c; din <= 32'h8a1eac09;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h044; din <= 32'h612d929e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d6; din <= 32'hf1991563;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08b; din <= 32'hf0ec106e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h173; din <= 32'hb8bf60d8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3fe; din <= 32'hf020e4cf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h276; din <= 32'hb8951f65;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h127; din <= 32'h5fe6cc36;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h32d; din <= 32'hb615c153;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0cc; din <= 32'hc3cf9b73;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h34c; din <= 32'hfb9e8027;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2dc; din <= 32'hfdc5a74e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h237; din <= 32'he7f6f589;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h36f; din <= 32'h512c259f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d5; din <= 32'hf8fce52e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h052; din <= 32'h00c25331;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00d; din <= 32'h08296aef;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h39f; din <= 32'hb514b895;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e6; din <= 32'h1a059a29;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h28b; din <= 32'h27c51153;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h11b; din <= 32'h256de08f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h318; din <= 32'h3ba48d31;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h174; din <= 32'h62958494;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3be; din <= 32'h7b8f155b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0fa; din <= 32'h776d23f1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h005; din <= 32'hd5cd7c3b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h076; din <= 32'h1d2d6ff9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h010; din <= 32'h52492cad;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h181; din <= 32'h4b876012;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b4; din <= 32'h0c59d4fc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ad; din <= 32'h01310cc8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h148; din <= 32'h2a5806d7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h25a; din <= 32'h34b02bf7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h125; din <= 32'h963e8c77;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h30d; din <= 32'hb392a808;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h021; din <= 32'haacbc382;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h158; din <= 32'h508d7e09;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h309; din <= 32'hf4fca41d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f8; din <= 32'h81d9ea40;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c1; din <= 32'h6b73f0dd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c0; din <= 32'h33df0cee;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ff; din <= 32'h9b23ec70;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h316; din <= 32'h24e918d9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c2; din <= 32'hc32938b4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h07d; din <= 32'h58995b58;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ef; din <= 32'hbb251893;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h300; din <= 32'h6528bee7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h025; din <= 32'h81fab18e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h34f; din <= 32'hca2177d6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h086; din <= 32'h64cd7c16;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h01b; din <= 32'h38cbd35a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h129; din <= 32'hbc008115;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h19d; din <= 32'h6244bdc2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h039; din <= 32'hdcffeba5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h065; din <= 32'h0c4bf2e6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d6; din <= 32'h14310b5a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c3; din <= 32'h64ba3216;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h120; din <= 32'he141cb1f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38c; din <= 32'haa6d5be6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ab; din <= 32'h456c10cd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h179; din <= 32'h1dcce36f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ec; din <= 32'he1522499;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h39c; din <= 32'hc216bca6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h103; din <= 32'h0fb6592b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h298; din <= 32'h05389e95;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38e; din <= 32'haf80146d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a9; din <= 32'h659ed1cd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h394; din <= 32'h9330c7cf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00c; din <= 32'hb1d6c43a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h334; din <= 32'hb700ec17;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h21c; din <= 32'h15e8ba6b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h222; din <= 32'h0346c86f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h335; din <= 32'hb309e0d6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h182; din <= 32'hec6dae37;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h311; din <= 32'h70a07169;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h183; din <= 32'h43845f81;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18a; din <= 32'h71f0bfe1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b9; din <= 32'ha043bc84;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h03a; din <= 32'hed7c975f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h359; din <= 32'h740cdadc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h104; din <= 32'h53fbad49;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e7; din <= 32'h151cc705;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h046; din <= 32'h7e27496f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h019; din <= 32'hdc7a6038;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c2; din <= 32'h1da0d3d4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23e; din <= 32'h158f03aa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08e; din <= 32'h9d813e53;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h33f; din <= 32'h7d0720de;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h26e; din <= 32'habfd7fd3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h33e; din <= 32'h636001ca;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0da; din <= 32'h1c2d22ee;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h359; din <= 32'hd42fa125;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h140; din <= 32'he8e9311f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ec; din <= 32'h22244eeb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d5; din <= 32'h3ad93c02;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h364; din <= 32'h59ef6acd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h002; din <= 32'h6410eaf5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1db; din <= 32'h219f3401;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38e; din <= 32'h00a51f09;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h344; din <= 32'h3dc45fbc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h077; din <= 32'hb13f709f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2a1; din <= 32'h74b3162c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h212; din <= 32'h81fa6eee;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h054; din <= 32'hac29b510;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18b; din <= 32'h9315ae0b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h02c; din <= 32'h45516ecd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h058; din <= 32'h15d43622;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f6; din <= 32'hca2a4d65;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37f; din <= 32'h9cf159c7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h368; din <= 32'h57127245;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e5; din <= 32'hd30a4145;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22f; din <= 32'h03b8d228;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b3; din <= 32'h896cd07f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f2; din <= 32'hd93739bb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h351; din <= 32'h224c5d6e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h048; din <= 32'h372925f3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ea; din <= 32'hb2d50057;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h358; din <= 32'hcad4b3d2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h10d; din <= 32'hd5450a19;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h287; din <= 32'h5a644a6f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h150; din <= 32'hcf3b67a9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c0; din <= 32'h2627c8ad;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h01d; din <= 32'hd1ffcdba;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h005; din <= 32'ha3db798d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d5; din <= 32'h6754fc12;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h13d; din <= 32'h6e786a9c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h288; din <= 32'h4147f99d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e3; din <= 32'h675aad10;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h197; din <= 32'h0715d2bc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d1; din <= 32'h3483ad9f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h35d; din <= 32'h1b479df7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h26f; din <= 32'h9862b9e3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h03e; din <= 32'hc6f41a50;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3cc; din <= 32'h2f800195;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h36a; din <= 32'heb256394;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h132; din <= 32'h5d264110;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h03c; din <= 32'hfb2c78d9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37d; din <= 32'h21d75ffa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h003; din <= 32'h71b20c94;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h330; din <= 32'hc1a630eb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b6; din <= 32'h733e670d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h206; din <= 32'h371d85b8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b6; din <= 32'h37fd2be8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h118; din <= 32'hee1f15a3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h15e; din <= 32'ha609f0e6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a3; din <= 32'h606bdeac;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e6; din <= 32'h9c7d0b7d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38d; din <= 32'ha3f1bf3d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h25a; din <= 32'h5d8fa91f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ad; din <= 32'h2c9386fa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h222; din <= 32'hebb1a8c8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h06e; din <= 32'he6ce5f3b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0fa; din <= 32'ha6c36d82;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h11c; din <= 32'hfda328ac;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a3; din <= 32'h3d4d4b50;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31c; din <= 32'hee83e112;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c7; din <= 32'h0e17795c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f2; din <= 32'h86900b43;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2bf; din <= 32'h8f226d01;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23a; din <= 32'hfc68a8bb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h25f; din <= 32'hd499e29d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h05b; din <= 32'h3fe9f06c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a5; din <= 32'heb70f9a6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c2; din <= 32'hb95dbd25;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3be; din <= 32'hee86ad5f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h076; din <= 32'h5ecd17de;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h29b; din <= 32'h94f0b657;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h286; din <= 32'h935de56a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h175; din <= 32'h7048a7c4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h029; din <= 32'hbeb18037;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16d; din <= 32'h255ac26f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h203; din <= 32'h8603332b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h036; din <= 32'h2fc0debf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22d; din <= 32'h07983fe4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h325; din <= 32'h290041d3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h34d; din <= 32'hc639a852;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h12a; din <= 32'h372c3c57;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ba; din <= 32'hfa5095c9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0dc; din <= 32'h824d3f39;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h269; din <= 32'h67f79e36;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h114; din <= 32'h67ed45ca;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h089; din <= 32'h4eb6ee28;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h323; din <= 32'h5b1c49c5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b1; din <= 32'h466790ea;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a3; din <= 32'h3da2124d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h07d; din <= 32'h9d8f9a5b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h108; din <= 32'h8c700765;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e8; din <= 32'h0d32049c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c3; din <= 32'h9f4154a9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h031; din <= 32'h85ef1386;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h306; din <= 32'hcaea2ab8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ed; din <= 32'hb31a7d94;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a6; din <= 32'h3cd95221;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e0; din <= 32'hdd2b7a5f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h153; din <= 32'h948e17a3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h097; din <= 32'h577177d5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h39d; din <= 32'h44e507d4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f9; din <= 32'h9ace50d7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h295; din <= 32'h6e2c2f0e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h337; din <= 32'h28c30df9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h256; din <= 32'hebd85a92;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h090; din <= 32'h82536902;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3fd; din <= 32'hc2a30cc8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a3; din <= 32'h34b361ea;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h243; din <= 32'h7e6eef51;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f7; din <= 32'h9442974d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h197; din <= 32'h844f0489;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h39c; din <= 32'hd5f9b465;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h216; din <= 32'h6a68fdd4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h366; din <= 32'h14c3ab00;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h05a; din <= 32'h2c158125;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h094; din <= 32'he74d342a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h213; din <= 32'haad06c49;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3aa; din <= 32'hf5682763;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0fd; din <= 32'hf0802f07;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h378; din <= 32'hd6ef8f4f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h277; din <= 32'h096b8efb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h06f; din <= 32'ha2ba9498;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h343; din <= 32'h00add296;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h35b; din <= 32'h5422f3e7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3dd; din <= 32'hefac0d52;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h092; din <= 32'h3d30c93d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c0; din <= 32'hf38fbc06;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c0; din <= 32'hea495be7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3cd; din <= 32'h32287a4e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h213; din <= 32'hcab40576;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0af; din <= 32'h850ee5a1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h092; din <= 32'h3b1ca09f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e7; din <= 32'h095e5a09;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c4; din <= 32'h0a6ad83d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h168; din <= 32'h6f2aab12;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d9; din <= 32'h0e956ee3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2a3; din <= 32'h25fc3b46;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h201; din <= 32'hca544311;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h25a; din <= 32'h0ad0ced8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2fb; din <= 32'hccb10733;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e8; din <= 32'hd07be8ff;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h367; din <= 32'h44a72e72;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h246; din <= 32'h4a261f34;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h19b; din <= 32'hff491f94;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h036; din <= 32'h5d72222d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h11c; din <= 32'h4278e9ae;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0bf; din <= 32'haea4ceb7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f2; din <= 32'h4123e268;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h265; din <= 32'h959541e4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h006; din <= 32'hf35fcc3b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h092; din <= 32'hd3d031a1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a1; din <= 32'h6f038d32;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08c; din <= 32'hc230fba1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b1; din <= 32'h931c7a14;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1fd; din <= 32'h5f24ac5e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h154; din <= 32'h1fe8aa60;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f4; din <= 32'he5b4e5a8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a0; din <= 32'h0a20cf1a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b3; din <= 32'hf2ace142;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ac; din <= 32'h1c4c4d75;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h29b; din <= 32'h14dffac0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h29c; din <= 32'he64b536b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h367; din <= 32'ha1e8ed11;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f0; din <= 32'h8f239161;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ae; din <= 32'h44aac95e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h231; din <= 32'hb0fbfb9c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b8; din <= 32'h8e0c2ba0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h175; din <= 32'h90e7040e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2a4; din <= 32'h44f57b2e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h004; din <= 32'he48ef68b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f7; din <= 32'h073ba634;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ec; din <= 32'hd8e74160;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e8; din <= 32'h7fc3359e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h35b; din <= 32'h7a69c2fe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h26f; din <= 32'h6304cd13;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ea; din <= 32'hf168fcee;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h201; din <= 32'hf02bc2be;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h297; din <= 32'h0b9f9531;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d6; din <= 32'hc77e221e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h265; din <= 32'h5fc1d447;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h292; din <= 32'he0559300;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h149; din <= 32'h5e2f3ac9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h174; din <= 32'h1053c0cd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h326; din <= 32'h63ec4d3e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h037; din <= 32'h6fac7972;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e2; din <= 32'h1b091ecc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h201; din <= 32'hbd07ec09;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f3; din <= 32'hfcd6197d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h32e; din <= 32'hf0bef327;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h34a; din <= 32'h67e88581;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b9; din <= 32'h3bbeba8d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d2; din <= 32'h0613a906;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e1; din <= 32'ha9668cd6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08c; din <= 32'hd031ae01;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h07b; din <= 32'hed81d53b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c1; din <= 32'ha0f92d7a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h037; din <= 32'hd1fb3fc7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b9; din <= 32'ha126f3d5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38f; din <= 32'h7b554b19;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h105; din <= 32'ha82ae254;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h314; din <= 32'h3faf4677;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h094; din <= 32'h1d562528;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h020; din <= 32'h65175187;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ac; din <= 32'h22a9b338;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h09e; din <= 32'h6cf79768;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a0; din <= 32'hb3cc30eb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b7; din <= 32'h3ced1f32;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h272; din <= 32'hfc6d71ca;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h036; din <= 32'h6731147d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h323; din <= 32'h9035c4ce;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h100; din <= 32'h1d6493bf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3fb; din <= 32'h98ee3d7f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h088; din <= 32'h054bd73c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f7; din <= 32'h55ee967e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h120; din <= 32'h168af9be;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h198; din <= 32'h3a1b3745;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h05f; din <= 32'hf73b7f7c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2a1; din <= 32'h04a77862;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h142; din <= 32'hdc706908;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h278; din <= 32'h9a07f1fa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37a; din <= 32'h0a1a435f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h13b; din <= 32'hd32397a6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b7; din <= 32'h03e8f065;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0bc; din <= 32'hd1bc640d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1cd; din <= 32'hf5b8ff1c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h04a; din <= 32'hc1d8075c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h163; din <= 32'h4af98060;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c1; din <= 32'hc468e724;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a1; din <= 32'hc20384d4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h338; din <= 32'h24d44c99;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1bd; din <= 32'h15a4ff66;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ab; din <= 32'h2b553f7a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h224; din <= 32'h846142b8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f3; din <= 32'hb69ca4ea;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h040; din <= 32'hd9437329;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a1; din <= 32'h58b4c9a5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2a7; din <= 32'h402ea5c7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e3; din <= 32'hbb94095f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h124; din <= 32'h1e8d18ce;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b7; din <= 32'h43dfa5fe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22e; din <= 32'hedc28e6d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h380; din <= 32'hf1450319;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h380; din <= 32'h6d005ca1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h34d; din <= 32'h5e95819f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c5; din <= 32'hc882382c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ff; din <= 32'hc1ba988c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22c; din <= 32'he651bfad;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h29f; din <= 32'hfa91605a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h015; din <= 32'h00639176;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3fc; din <= 32'h4fce61e9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h29d; din <= 32'h7fd28d42;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h397; din <= 32'h0944f1fc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h145; din <= 32'he6c04fb5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h20f; din <= 32'ha87c222a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b9; din <= 32'h49e1392a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h19a; din <= 32'hb603f7b8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h069; din <= 32'h4da793e5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h019; din <= 32'h4b06b753;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1be; din <= 32'hd5641499;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h372; din <= 32'haa7195be;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3fb; din <= 32'heff49d00;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h398; din <= 32'h2c5ddfe2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2a2; din <= 32'h390dd9f2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h369; din <= 32'h518544a3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h32a; din <= 32'he00fa189;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e1; din <= 32'hef9f8793;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h267; din <= 32'h616cd96a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h264; din <= 32'h6b1442ba;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h382; din <= 32'h0c009d07;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h377; din <= 32'hbd821d63;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h210; din <= 32'h44d01183;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h01c; din <= 32'h61fe3fe5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h360; din <= 32'h8dec60e2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h04d; din <= 32'h1921843d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00b; din <= 32'hf634cfae;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ef; din <= 32'hbd4c210d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h379; din <= 32'h226ddbaa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h12d; din <= 32'hf3c7cc31;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h245; din <= 32'h316e3c78;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b2; din <= 32'hea77c90c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h251; din <= 32'h3f6b7bf5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h012; din <= 32'h5cc1a833;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a2; din <= 32'h235ae2c1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f8; din <= 32'h05b99131;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b7; din <= 32'h42376c14;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d5; din <= 32'h3f7d5ea9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h362; din <= 32'ha4e0df40;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e9; din <= 32'hcb434348;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c0; din <= 32'h1d487389;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h005; din <= 32'h4cd9d17f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h103; din <= 32'h94cffb2d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c5; din <= 32'hc3b339ad;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ad; din <= 32'hb67c7cee;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b3; din <= 32'h881bb84c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h05f; din <= 32'h6e674d67;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h208; din <= 32'h7c393de1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h01c; din <= 32'haefa483b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ed; din <= 32'h87bec025;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h06b; din <= 32'h43338138;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h332; din <= 32'hd489ec79;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h280; din <= 32'h9ae17ca7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d5; din <= 32'h29b5d94b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h353; din <= 32'h89ff0e3c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h219; din <= 32'hd0db697e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3de; din <= 32'h0948690a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d2; din <= 32'h2917e1cf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c4; din <= 32'h8f4afe6b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h246; din <= 32'h0472d159;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h312; din <= 32'hc501de7e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h321; din <= 32'hbde6cd7f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a1; din <= 32'hed0d4e9a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f3; din <= 32'hed127349;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00d; din <= 32'h8392c118;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h059; din <= 32'h0833ab79;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f4; din <= 32'h0809b121;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h184; din <= 32'h0d170f85;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c0; din <= 32'hfdcf0797;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h247; din <= 32'h16a7ccbd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2fe; din <= 32'hb58cad4f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ec; din <= 32'h58aeef32;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b7; din <= 32'h8243efc8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31b; din <= 32'h2e979887;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h207; din <= 32'h74c4023e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h138; din <= 32'hb2753f65;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h28e; din <= 32'he2c90ed6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h022; din <= 32'h4248b7a6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h14c; din <= 32'h95be02a1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h12b; din <= 32'h76c98e7d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ec; din <= 32'h53e6a402;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h19a; din <= 32'h931d3c86;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h07c; din <= 32'hdf36c32d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h165; din <= 32'h4615115b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h35d; din <= 32'h275e3d2b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a5; din <= 32'hb2324f09;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h01e; din <= 32'h7e2c6cfe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18a; din <= 32'h6e0d4237;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h211; din <= 32'h3f26edb7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c0; din <= 32'h1d39fd2a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h133; din <= 32'hdce85c71;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1cf; din <= 32'haa9e11f4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h064; din <= 32'h1df913b7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h33f; din <= 32'hdeb81f45;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b9; din <= 32'h2913291f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h191; din <= 32'h067c3101;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3de; din <= 32'h91c49b8e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h090; din <= 32'h2f03029a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h04f; din <= 32'he2d5d13d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h231; din <= 32'h272c75d6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h29d; din <= 32'hc0a113c4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h160; din <= 32'h55539e42;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2a2; din <= 32'h2b9c91fa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h341; din <= 32'h95637c7f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2df; din <= 32'h10cfdb0d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2dd; din <= 32'h633cba05;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08a; din <= 32'h40491e10;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h02a; din <= 32'hcd04c545;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h33c; din <= 32'h76fcfa02;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h193; din <= 32'h653eda45;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h04e; din <= 32'h6effcc9f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h038; din <= 32'hd42ef739;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h24f; din <= 32'h8bf8504c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h04d; din <= 32'he2a98a86;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h06e; din <= 32'hcfbd9e9d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h293; din <= 32'hc900c3a9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ef; din <= 32'h89c880ea;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h109; din <= 32'h805361fe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ea; din <= 32'h3f292be9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h28e; din <= 32'h628300bb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2cf; din <= 32'h4c558616;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h13f; din <= 32'h068f7b2c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h067; din <= 32'h624cfe6e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31d; din <= 32'h1996b409;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h03b; din <= 32'h2f28f28d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h124; din <= 32'hc4e69b6d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h095; din <= 32'h01188aca;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h167; din <= 32'h298faf0e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h32f; din <= 32'h5e3c3610;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h069; din <= 32'h2d73cb24;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b9; din <= 32'h3c643b12;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3cb; din <= 32'hf9adf3f5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2eb; din <= 32'h0239a9d0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h156; din <= 32'h2052381c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ac; din <= 32'h423bab4f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h07b; din <= 32'h27b0236c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h167; din <= 32'ha24fd81c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c4; din <= 32'hec40fa8c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23d; din <= 32'h86a3e5a9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h17b; din <= 32'hc5bf6716;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h127; din <= 32'hfc3661de;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h097; din <= 32'he84996f8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a9; din <= 32'h194bc5a4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b8; din <= 32'h8f6016d0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d3; din <= 32'h9029c31a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ff; din <= 32'hdc11b511;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00c; din <= 32'h4f2d9910;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h359; din <= 32'h2315d8c9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h143; din <= 32'h56796489;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f4; din <= 32'h8e42be77;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0cc; din <= 32'hb32718b4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h305; din <= 32'hc3a6f493;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h13c; din <= 32'h42222fc2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2bb; din <= 32'h17e1db16;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h319; din <= 32'h7920db71;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h221; din <= 32'hc193b1eb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h30a; din <= 32'h932754ba;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h162; din <= 32'h3483fcf4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a7; din <= 32'h744c725b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h132; din <= 32'hf3ea7b65;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c2; din <= 32'h40351609;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a6; din <= 32'hecd8eafe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h194; din <= 32'h50cbf827;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h313; din <= 32'h6fe1ab01;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18e; din <= 32'hdb188d55;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h371; din <= 32'h3c303705;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b9; din <= 32'h9d214ccd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h03c; din <= 32'h8e8d651e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h21f; din <= 32'h35b20770;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h021; din <= 32'hfdba54b3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e9; din <= 32'h56f88a2b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0eb; din <= 32'h7b5d303f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h008; din <= 32'hc87152d4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h237; din <= 32'h8e5c4c26;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ca; din <= 32'h4801cbeb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h056; din <= 32'h38ef32db;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h05e; din <= 32'hd0eca183;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h270; din <= 32'hb26b8472;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3cc; din <= 32'h243dbaf7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d0; din <= 32'h40c7bddd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h150; din <= 32'h705ac686;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h127; din <= 32'h8412b469;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h250; din <= 32'h95cc8969;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h200; din <= 32'h9546c4b7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h347; din <= 32'hdcbb57a0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h167; din <= 32'hb1994686;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h01a; din <= 32'hbb85b349;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h02a; din <= 32'h824fba9b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h01f; din <= 32'hd1f3187a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h26e; din <= 32'h7f798cf0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h352; din <= 32'he8fa5436;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h09f; din <= 32'hd0d8938c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0cf; din <= 32'h6fcbbc92;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h36a; din <= 32'h934f1953;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h199; din <= 32'h7484a06a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h06c; din <= 32'h3c1d202d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a1; din <= 32'hf319df2e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h253; din <= 32'hedf5dc43;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b3; din <= 32'h77a509f1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h113; din <= 32'h29cc2c2f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c6; din <= 32'h31b73576;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h13f; din <= 32'hd2153ca7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h24d; din <= 32'h120ddbae;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f3; din <= 32'h79caf501;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h193; din <= 32'hfa7602f3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f7; din <= 32'hbb396bf6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h27c; din <= 32'h7115029a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h390; din <= 32'h59f98308;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0da; din <= 32'hb87e64f6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h191; din <= 32'ha6e7133b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h124; din <= 32'hcd8ec16c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ee; din <= 32'hb95130b4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ba; din <= 32'ha6de2689;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0fb; din <= 32'h2298f06b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b9; din <= 32'h3036aa26;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h34f; din <= 32'hf59896ff;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00f; din <= 32'h82449197;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08a; din <= 32'h5aa46aa5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h25b; din <= 32'h6dc2abf9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08b; din <= 32'h466ff574;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h084; din <= 32'h6201095f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h235; din <= 32'h2cfc1afd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h225; din <= 32'h54c4faaa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h24e; din <= 32'h91f25a3a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a0; din <= 32'h117fe702;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h09d; din <= 32'hbf3d38df;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37f; din <= 32'h89b11e85;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f0; din <= 32'h64d5a1ac;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f7; din <= 32'h11fa2a2c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f4; din <= 32'h202713cb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h320; din <= 32'h3128906c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h26d; din <= 32'h49f42460;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h35e; din <= 32'h64c3ff8d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ba; din <= 32'h53d1123d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e3; din <= 32'hf121e203;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h33e; din <= 32'hea496fb1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h028; din <= 32'hab2b0596;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d6; din <= 32'hdf6d47e0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h135; din <= 32'h5e8efd17;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c1; din <= 32'h312e4c3c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a3; din <= 32'hfa1aaf3b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0cf; din <= 32'h8cca9dcb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h089; din <= 32'h4b2c4dd3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h33e; din <= 32'hcb95f5cd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h318; din <= 32'h3d8f580d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h165; din <= 32'ha039c34f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23e; din <= 32'h02ecf373;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e9; din <= 32'h669bc81c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a3; din <= 32'h5c0c96e6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h007; din <= 32'hf40b817c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h322; din <= 32'hb6b1d1b4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e3; din <= 32'hc742e3d2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b1; din <= 32'h8bb6b5b7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h386; din <= 32'h51904839;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h07b; din <= 32'hf2f9eff6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h399; din <= 32'h09c8c730;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h215; din <= 32'he53bbd42;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a4; din <= 32'h9012cbfa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h335; din <= 32'hd89ff0fc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h049; din <= 32'haec7db87;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h069; din <= 32'h6c08cf32;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h277; din <= 32'h602f09ed;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h300; din <= 32'h435d10ef;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00e; din <= 32'h27f56b4a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h27c; din <= 32'h0a861a25;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d0; din <= 32'h1bff5a95;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23e; din <= 32'hf0f18c12;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f1; din <= 32'h800be33e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h212; din <= 32'h4f38bee6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e2; din <= 32'h5bb3df0e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e5; din <= 32'h3d4a7baa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h282; din <= 32'h3b2782cb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f4; din <= 32'h2aec82d4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c2; din <= 32'h639f2637;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e1; din <= 32'h630fad82;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h043; din <= 32'h31f72c96;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h353; din <= 32'h04b11765;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h370; din <= 32'ha8794f8f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h357; din <= 32'hb4318d60;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h034; din <= 32'h6316bcfd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b8; din <= 32'hcfe7e9a1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16b; din <= 32'haf387e43;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h338; din <= 32'h9332c52e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2af; din <= 32'h94324692;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h321; din <= 32'h5ac22a07;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h334; din <= 32'h42a3bbc7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h062; din <= 32'h2617b108;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d3; din <= 32'he58853e6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h124; din <= 32'h09722609;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h02b; din <= 32'hc12d6151;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0fd; din <= 32'h9e3edc1b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h126; din <= 32'hc8550691;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h27f; din <= 32'hb282e932;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h095; din <= 32'h98a323df;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h232; din <= 32'h0834fe22;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h217; din <= 32'ha6b3d017;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h138; din <= 32'hc9562ee2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23a; din <= 32'h1eca8983;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18c; din <= 32'h426f3341;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2af; din <= 32'h11822e8b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3cb; din <= 32'h60990aaf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d1; din <= 32'hbe91deb1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h162; din <= 32'hf2b050d8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ee; din <= 32'h6083722f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h279; din <= 32'h6ff6fc01;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c9; din <= 32'h23862a03;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h224; din <= 32'hb38fc521;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h21a; din <= 32'h0dcec027;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h181; din <= 32'h36f3b9b6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3be; din <= 32'haf8303d0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h257; din <= 32'h8a7056f3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18b; din <= 32'hdc5195e6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31a; din <= 32'h81923277;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d1; din <= 32'h7f609ac3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b0; din <= 32'h172a655a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22c; din <= 32'h038ffcc2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h27a; din <= 32'h4570614c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ef; din <= 32'h591ae363;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a7; din <= 32'hb6ce4cea;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ef; din <= 32'hdea068e7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h01e; din <= 32'h232e63bb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h150; din <= 32'h1be08b87;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h279; din <= 32'h6bfdfbde;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h03e; din <= 32'hcbea8225;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h122; din <= 32'h4372393b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h27e; din <= 32'hbb81342f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0dd; din <= 32'h1363e048;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3fa; din <= 32'hb8a676a3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h06f; din <= 32'hf87aee1a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h090; din <= 32'h32319fa2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h134; din <= 32'h1e08f0a5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ee; din <= 32'h61b89a30;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h205; din <= 32'h2621de75;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h210; din <= 32'h9e570756;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38a; din <= 32'h0b80f634;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h253; din <= 32'h6d8f22e9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h190; din <= 32'hd8b02d61;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h318; din <= 32'h75711f83;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a6; din <= 32'hc800c84f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b4; din <= 32'h02d5eb3b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e8; din <= 32'he0222251;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h363; din <= 32'h31de6650;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1da; din <= 32'h983cfb53;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1fd; din <= 32'hba09d811;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31e; din <= 32'h0c6e265b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h300; din <= 32'hbe936b34;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h073; din <= 32'hf87729af;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h005; din <= 32'h58c2c53e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h201; din <= 32'h3d3d021f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37c; din <= 32'hedc8656f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22e; din <= 32'h9b259dbd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h344; din <= 32'h614fc61f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h19f; din <= 32'h9af9a32c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h229; din <= 32'hce7a5431;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c3; din <= 32'ha051ddff;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c9; din <= 32'he26f2e3d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h05b; din <= 32'h3b84dd74;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08e; din <= 32'h3312fb10;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3cf; din <= 32'h7b004db8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h115; din <= 32'haf17d097;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0cf; din <= 32'hc4d963e6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h270; din <= 32'h9070f2f3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h369; din <= 32'h5e2aa523;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h07d; din <= 32'hc423fcf4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a1; din <= 32'h5055db35;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h293; din <= 32'h30d2d346;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h03c; din <= 32'hd7df0c3a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h018; din <= 32'h7a0c73e3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f6; din <= 32'h4ced24b3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f3; din <= 32'h433141d7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0bf; din <= 32'hc8b612eb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d4; din <= 32'hffae3250;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ff; din <= 32'hd7e99a75;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a5; din <= 32'h59592d59;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00b; din <= 32'hce73988b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18f; din <= 32'h9e4041f7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h39e; din <= 32'hf026f2b7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ee; din <= 32'hb16fe346;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d5; din <= 32'h2d26f570;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h367; din <= 32'h2dbcd3d3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h172; din <= 32'h67624827;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h14c; din <= 32'h2f2ee6bf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f2; din <= 32'h438ec783;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h07e; din <= 32'h4ec8ec66;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a0; din <= 32'ha76250a6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h01f; din <= 32'hadbc8275;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a7; din <= 32'h6d4c65bd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h267; din <= 32'h4bdcd9ca;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1dc; din <= 32'ha5aa2bcc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h01a; din <= 32'h62427f50;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1cf; din <= 32'he15b9396;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h09b; din <= 32'heda4e0f6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h018; din <= 32'hb06c9107;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a0; din <= 32'hea360aeb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h181; din <= 32'h8b3852a6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h30f; din <= 32'h5c52f44b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2cf; din <= 32'h2717cb21;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h34c; din <= 32'he814371c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h13a; din <= 32'h73f8cf10;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d7; din <= 32'hf9d3048c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d7; din <= 32'ha532507a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h184; din <= 32'h96cad787;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h374; din <= 32'h5e16ed41;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h091; din <= 32'he3c96d15;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c7; din <= 32'hc9a331d6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h205; din <= 32'h3684ecd3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1fb; din <= 32'h869f4164;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h01f; din <= 32'he118edc7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h151; din <= 32'hea5602e7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a9; din <= 32'hdfc26593;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a9; din <= 32'he8c81b95;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0de; din <= 32'h7295ba6f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h041; din <= 32'h5987d736;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h17a; din <= 32'haec2e8d6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c2; din <= 32'hc05af7fa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h143; din <= 32'h0dc8b3b0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f6; din <= 32'h3b6b74d6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h26d; din <= 32'h1ae4aaf8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h200; din <= 32'h4fd17bd0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h28b; din <= 32'h9c0426a8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h325; din <= 32'h7df62000;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h33d; din <= 32'h6743e5cf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0eb; din <= 32'ha55f0001;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a3; din <= 32'h80d58423;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h19c; din <= 32'h6f240950;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h33f; din <= 32'hff338322;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h002; din <= 32'h36701d8f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1cc; din <= 32'h22d8569d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h103; din <= 32'h7958ead1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h24e; din <= 32'ha7142853;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h03b; din <= 32'hfa09d30c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f3; din <= 32'h096d018a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e4; din <= 32'hd4c2da63;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h083; din <= 32'hec2e943a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3bb; din <= 32'h2c35f53f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d7; din <= 32'hdab80d62;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3bd; din <= 32'h7b478dd3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h009; din <= 32'hf5ef9b3b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h356; din <= 32'h1edff798;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h061; din <= 32'h8e31aca9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h079; din <= 32'h1dad8a75;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h133; din <= 32'hbbbd67fe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a4; din <= 32'hf7c9d36c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h246; din <= 32'h03e0193c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b4; din <= 32'h359c4e59;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h06b; din <= 32'h4bb83227;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b0; din <= 32'hfeab69a4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h30d; din <= 32'h4c9d6a7c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ea; din <= 32'h89a09455;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h19f; din <= 32'h1206ea9f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h253; din <= 32'hf8327f32;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c1; din <= 32'h71d77ea3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h06e; din <= 32'ha905c752;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h11d; din <= 32'h3c168dbd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0cc; din <= 32'ha40043b6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2fe; din <= 32'h48050a50;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h13a; din <= 32'h4939145b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h009; din <= 32'hfd020afa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h317; din <= 32'h8c327ef9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1fd; din <= 32'h4a2c1c95;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31b; din <= 32'h819de2fe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h09f; din <= 32'h81ffaef5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c2; din <= 32'hf32bba31;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d1; din <= 32'he06c7568;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h219; din <= 32'hb2771472;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h061; din <= 32'h344ddad0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h399; din <= 32'h6b5698b3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38f; din <= 32'h14f53412;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h17d; din <= 32'h7b9d547f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c5; din <= 32'hb68f75f7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c0; din <= 32'he2852b18;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2aa; din <= 32'he303d743;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0fa; din <= 32'hc5f3366d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e7; din <= 32'hf4ceb8a6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h111; din <= 32'h023f56f3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h027; din <= 32'hf2a51be6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h335; din <= 32'hf151d450;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h193; din <= 32'h5aeb2272;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d7; din <= 32'h3dde7a95;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16b; din <= 32'h37498447;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h391; din <= 32'h3299eee1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a0; din <= 32'hc2dd6e90;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00d; din <= 32'h5441f2c2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h348; din <= 32'h0f787977;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h111; din <= 32'hd06def27;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3bd; din <= 32'hb80d14d8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h183; din <= 32'hb56ebf9f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h014; din <= 32'hbd1f5d41;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d9; din <= 32'h95a6c475;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2a4; din <= 32'hea5ab3a7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h195; din <= 32'h6162a80d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h212; din <= 32'hbb2065e0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18d; din <= 32'hc40e5e01;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h159; din <= 32'h84653ff2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h201; din <= 32'hd54e2e8c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a9; din <= 32'h6a57af1f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e4; din <= 32'h54faa357;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h229; din <= 32'hc37ba716;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h196; din <= 32'hb9845599;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h25b; din <= 32'hdf979f73;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e7; din <= 32'h6aadeb62;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c6; din <= 32'hb906c837;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08b; din <= 32'h343e7b2c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h286; din <= 32'ha496692b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h20c; din <= 32'h7e96acc7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0eb; din <= 32'h27365d57;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16d; din <= 32'hac278fac;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d0; din <= 32'h0d334484;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h36b; din <= 32'h980c21b6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h238; din <= 32'h078186b2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h240; din <= 32'hc0474cec;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h224; din <= 32'h91607699;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e5; din <= 32'hd4f4dd23;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a0; din <= 32'h03ccd76f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3df; din <= 32'hb1536841;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h018; din <= 32'h0b979c7e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ba; din <= 32'hba65be78;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1bb; din <= 32'h42146e92;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h211; din <= 32'h93f15fb0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h283; din <= 32'h5a6e1b38;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08f; din <= 32'h083853ed;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h296; din <= 32'h5d144d05;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f4; din <= 32'h17092898;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d0; din <= 32'hc1c5e8d2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ee; din <= 32'hc2c54916;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c0; din <= 32'ha6cc4b83;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h242; din <= 32'h1010788c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ca; din <= 32'h4c1f0c9a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3bc; din <= 32'hd103201a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3eb; din <= 32'h6c146655;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00f; din <= 32'h9d83d152;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ed; din <= 32'hf30743a9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h003; din <= 32'h5bcc614d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h34c; din <= 32'h30de3d67;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0fc; din <= 32'h48f63df8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h11b; din <= 32'hbe9cb5a4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h166; din <= 32'hfdc8472a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ba; din <= 32'h4da2bd2b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31d; din <= 32'hd8d20ba6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h272; din <= 32'ha7556d5f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h35a; din <= 32'h1d6dd004;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h238; din <= 32'h23e1ce65;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ce; din <= 32'h6c16e6be;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d2; din <= 32'h2184988e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h031; din <= 32'hdb15524a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h280; din <= 32'ha2d9ac79;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h09b; din <= 32'h785165f6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2dc; din <= 32'h9c38abf7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h14e; din <= 32'h06b486b4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h11e; din <= 32'hafc491bc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h055; din <= 32'h666bf0e9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h266; din <= 32'h12abf778;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h079; din <= 32'h7f27ddc7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h110; din <= 32'h8a1e3767;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0cd; din <= 32'h31255037;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h215; din <= 32'h61fa47b8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e6; din <= 32'h3863a336;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h136; din <= 32'h6942f687;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b7; din <= 32'h5e73d3c9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f6; din <= 32'ha9714f3b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h218; din <= 32'h3c432937;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h000; din <= 32'hd847944e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h296; din <= 32'hc3b9a8aa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h167; din <= 32'he8b5810a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f5; din <= 32'h2a5ac39e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h178; din <= 32'h7556768b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d4; din <= 32'h083e8acf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0fd; din <= 32'hd126e5db;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h01d; din <= 32'h2cfe033c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h014; din <= 32'h5a25b3e5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h24b; din <= 32'h7ff047e2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h075; din <= 32'heb7b9b7d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0db; din <= 32'hb7a7a4c9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h36e; din <= 32'hebcc4e10;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h006; din <= 32'h3dff5926;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h263; din <= 32'h275d3b79;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h081; din <= 32'h17920394;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h088; din <= 32'hd8643802;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18b; din <= 32'h34e544ae;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h390; din <= 32'h82e75086;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h257; din <= 32'h5eee7695;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h003; din <= 32'hf6a61fe8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16d; din <= 32'ha5dff7fc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h019; din <= 32'h6937b7f7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h28d; din <= 32'h71723b9d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ee; din <= 32'h15b3809b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h171; din <= 32'h6ba515fa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h12f; din <= 32'h3a607c0c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h120; din <= 32'hfea000d3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22d; din <= 32'hc7cd6b42;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22b; din <= 32'h28481fbb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08c; din <= 32'h917d6c87;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h21b; din <= 32'ha24df1df;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a1; din <= 32'h9aea4997;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h323; din <= 32'h20b234bc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h178; din <= 32'h2ab2c4da;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h36c; din <= 32'h215839b1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0bd; din <= 32'h3863b722;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c2; din <= 32'h2e303d2f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c1; din <= 32'h2bedd882;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h19e; din <= 32'h028f68a4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h17c; din <= 32'ha0006f56;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h30e; din <= 32'h3b9af397;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a8; din <= 32'ha295d8f0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e1; din <= 32'hc07ab1ca;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h077; din <= 32'hc8016c9d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ed; din <= 32'h2fbf56cc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d4; din <= 32'h52f8e837;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h27b; din <= 32'h88e7f9d6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f9; din <= 32'h40617944;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h171; din <= 32'h527ad99d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h170; din <= 32'h74bc2b20;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h25d; din <= 32'h3daee8d0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h390; din <= 32'h6da4fdeb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ba; din <= 32'he5444975;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h189; din <= 32'hf9686859;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e6; din <= 32'h5fe8e1bd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h114; din <= 32'h5a58693f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d9; din <= 32'h646e1359;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08f; din <= 32'h43a5d120;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h160; din <= 32'hb5cf844f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h05c; din <= 32'hcadb27a5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h008; din <= 32'hbfb0cce5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b0; din <= 32'haacf0b0f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h341; din <= 32'hdc470e8e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h39b; din <= 32'hd171629b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h369; din <= 32'h47aa3ee2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h004; din <= 32'h6fd74614;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d2; din <= 32'h3ba36b27;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h071; din <= 32'h846d89a8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h214; din <= 32'h3e1920d5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h148; din <= 32'h029a48f5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h199; din <= 32'h9798ffcd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h234; din <= 32'h69176d3e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h185; din <= 32'h11601d3e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f1; din <= 32'hd812b3a0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h375; din <= 32'h1214d5d1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h131; din <= 32'hfa7cbe54;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h042; din <= 32'h7ac470e8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h273; din <= 32'h35cd12b0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a6; din <= 32'h50bead17;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h04a; din <= 32'h278f21c8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h138; din <= 32'h87fd3f51;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h205; din <= 32'hbd1625ec;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f5; din <= 32'h9959e709;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ba; din <= 32'habcdaad9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h222; din <= 32'hf0e6a203;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b2; din <= 32'h085a3049;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h089; din <= 32'h0c2f5ac3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b8; din <= 32'h748f4662;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h049; din <= 32'hff62e7b8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h01a; din <= 32'h3c3c5cdd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2dc; din <= 32'hd5a50910;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h397; din <= 32'h49f4307a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a4; din <= 32'h06279d77;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h26d; din <= 32'hc455225a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b5; din <= 32'hdd0281f7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h056; din <= 32'h929a9dfa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h341; din <= 32'had6a6105;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b7; din <= 32'hd861e3e2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h120; din <= 32'hb4b7270b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h11e; din <= 32'h005edf48;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h02b; din <= 32'h097b5a87;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ac; din <= 32'hff9f399d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h323; din <= 32'h4d492a9d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h395; din <= 32'h559b5280;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h178; din <= 32'h2804510e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h27e; din <= 32'hcd7991fd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h313; din <= 32'h69fb7035;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f8; din <= 32'h48e24c6e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h34e; din <= 32'h37551aa7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h34f; din <= 32'ha8b847a3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b8; din <= 32'h709cff5e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e0; din <= 32'hb14a1730;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3fc; din <= 32'h237296c4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h290; din <= 32'h261b5d1d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h02f; din <= 32'h4533bbf9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h270; din <= 32'h9d3444f8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h213; din <= 32'h8e390511;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h364; din <= 32'ha65d3469;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h352; din <= 32'hf7451345;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ad; din <= 32'h71d9d64b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h13b; din <= 32'h30d42277;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h13d; din <= 32'h8f858184;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37f; din <= 32'h90d698b9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h259; din <= 32'hf314e0f3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23b; din <= 32'h50310da8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h196; din <= 32'h498109fa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c9; din <= 32'hb4cf1b04;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h07e; din <= 32'h2abeac0c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3df; din <= 32'h4b9accc5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h083; din <= 32'h88c1ae26;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h009; din <= 32'h88488bdf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h391; din <= 32'h0c0bae1a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h088; din <= 32'h90dbc0c8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e0; din <= 32'h80eb05f9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0fc; din <= 32'h9ad75651;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b1; din <= 32'h24c348a6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h008; din <= 32'h69fc6f63;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h247; din <= 32'had693d9a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h35d; din <= 32'hdc65ada3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e8; din <= 32'hce5ce77c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h21e; din <= 32'h17e8a75f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00d; din <= 32'h7adf80db;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a8; din <= 32'h608e1a1c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e7; din <= 32'h12110037;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b1; din <= 32'hf850a6d4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b3; din <= 32'h940029a8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08a; din <= 32'hed3a263e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h103; din <= 32'h29e9cd06;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b5; din <= 32'h806b1def;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h036; din <= 32'he026bf3b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b0; din <= 32'hee345056;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ce; din <= 32'h59eb8874;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h245; din <= 32'h20d83084;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f7; din <= 32'h4ada1632;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h141; din <= 32'hef92b12a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0da; din <= 32'hbdd61726;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ea; din <= 32'hba7e0d6f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h204; din <= 32'hca230460;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2af; din <= 32'h7ad0e7f9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h14b; din <= 32'hf20dd137;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h376; din <= 32'h338afb80;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38f; din <= 32'h4e973e85;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a2; din <= 32'h0e5ab09a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3db; din <= 32'h1f179636;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ba; din <= 32'hf57cfec2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h072; din <= 32'h8aa444d5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1fa; din <= 32'h92fc44b1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h130; din <= 32'h34fdd534;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h355; din <= 32'h3766a729;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b1; din <= 32'he623a712;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b5; din <= 32'h5a3373b8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1db; din <= 32'h79634746;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c1; din <= 32'hc2579ddb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b1; din <= 32'h36b20579;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h315; din <= 32'hbac11481;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16f; din <= 32'h6741d4d2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h001; din <= 32'hf20649ee;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h33c; din <= 32'hd8ed0866;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h073; din <= 32'he43d4b46;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e2; din <= 32'h78399dc1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ec; din <= 32'hadf341f4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h033; din <= 32'h600d79a6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2a4; din <= 32'hee9d1d92;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h224; din <= 32'h57735009;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h306; din <= 32'h00f62c2b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3dc; din <= 32'h06d89810;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h294; din <= 32'h6507ccf3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16a; din <= 32'he60d3d85;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h284; din <= 32'he0752d63;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0fb; din <= 32'h49752ff6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0bf; din <= 32'h4952d0c7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c1; din <= 32'he587195b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h126; din <= 32'hf58ab6f7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h295; din <= 32'h891e65dc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3eb; din <= 32'h1f98a88b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38a; din <= 32'hc88bc91a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ef; din <= 32'hc31b45c3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h29c; din <= 32'h71c115fd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h169; din <= 32'h0c2bc48c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f9; din <= 32'hd58fabba;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h249; din <= 32'h516c002a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b1; din <= 32'ha64eb8b0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h340; din <= 32'h711cb5cf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h374; din <= 32'he8c18660;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h243; din <= 32'h57be24d7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h068; din <= 32'hd0760783;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h149; din <= 32'h16b42bf3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h198; din <= 32'hc3dfe97d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1dc; din <= 32'he1376c9c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1aa; din <= 32'h4f0ee615;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37c; din <= 32'h4ce9ddd3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ae; din <= 32'h81475046;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31e; din <= 32'haee9e225;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h25b; din <= 32'heb970e5a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37e; din <= 32'ha369d6d7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ae; din <= 32'hb251f18c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2a0; din <= 32'hac0191e0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d9; din <= 32'h3d4a7316;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h332; din <= 32'h19555f6b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h24b; din <= 32'h47940063;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h045; din <= 32'h0af67600;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1bf; din <= 32'h397ba51a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h251; din <= 32'h008ecd78;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00b; din <= 32'ha68dcc72;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h30f; din <= 32'h21a8f595;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h308; din <= 32'hd4366faf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h28d; din <= 32'h2af5ab59;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h003; din <= 32'h65b83a75;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h104; din <= 32'hde81f9ee;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b9; din <= 32'h655ac91b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b9; din <= 32'hc4624d91;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h15e; din <= 32'h92fae8c9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ba; din <= 32'hc28c93a4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h023; din <= 32'hed05e0df;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h057; din <= 32'h19132393;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h357; din <= 32'h08c99063;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h140; din <= 32'h781590c2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h291; din <= 32'h1a785810;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h221; din <= 32'h52884399;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b2; din <= 32'h610aaf79;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h131; din <= 32'h674fe4b1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0bc; din <= 32'hea56e565;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h243; din <= 32'h318ad70c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h258; din <= 32'h80b16999;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a7; din <= 32'h5f8250a7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38f; din <= 32'h8a9d4997;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ed; din <= 32'hc347e62d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h184; din <= 32'h244641a1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h236; din <= 32'hac4bcf1c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h388; din <= 32'h47c6229b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ae; din <= 32'hebff8b92;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h34f; din <= 32'h8f82f6a7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h208; din <= 32'hd4e771b0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h373; din <= 32'h8529824d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h224; din <= 32'hf4ce1be7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18e; din <= 32'h16b77d1b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h173; din <= 32'h74e5240b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b0; din <= 32'ha46cf800;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h117; din <= 32'hbed940f5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h124; din <= 32'h53e3f066;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3de; din <= 32'h6fb357df;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2a3; din <= 32'h22cd4a6f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c8; din <= 32'h00277bb7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h310; din <= 32'h45b428a4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h149; din <= 32'h283c6828;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h136; din <= 32'h8c7574de;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h236; din <= 32'h92b2c7c5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h388; din <= 32'h6f40ef44;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h149; din <= 32'h959f600c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0de; din <= 32'hbd613ae9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23a; din <= 32'h19af5237;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h191; din <= 32'hc6e5db4b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c8; din <= 32'h666ee9f2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h30b; din <= 32'h27768cb2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a7; din <= 32'hb1c7fe80;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b7; din <= 32'h71b51d83;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ba; din <= 32'h1be2e154;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h387; din <= 32'h50e7e211;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00d; din <= 32'h6facc7cd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h36f; din <= 32'hcc505349;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2fb; din <= 32'h1e8c9f3a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1fb; din <= 32'hafa4e6df;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h33a; din <= 32'h7c6ea535;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h394; din <= 32'h3c7bab67;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h293; din <= 32'hbf14b2c2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0dc; din <= 32'h17076a11;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h04b; din <= 32'h3901029a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08e; din <= 32'h46c9b971;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2de; din <= 32'hd922ad4b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f9; din <= 32'hc653804f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1bc; din <= 32'hfcceb13e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h35e; din <= 32'hd2073de1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h293; din <= 32'hbb225115;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f0; din <= 32'h327fa502;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3db; din <= 32'ha5aa5d67;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c1; din <= 32'h4bba8f87;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h13e; din <= 32'h0a3530a6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h32b; din <= 32'h254fca11;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h338; din <= 32'h40e1bd33;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18d; din <= 32'hbb289c00;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h25b; din <= 32'h630fceb1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f9; din <= 32'hcd5ce599;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h080; din <= 32'h479e2bcd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h01d; din <= 32'h952d5635;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h309; din <= 32'hbfb67d87;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a1; din <= 32'hf5acd0cf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b2; din <= 32'hdabde7d9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e7; din <= 32'he94201f2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h028; din <= 32'h7525c891;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h11f; din <= 32'hde462c24;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h098; din <= 32'h837ad77a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h218; din <= 32'hf6d02b31;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h218; din <= 32'h0c0dfccc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h066; din <= 32'hddb92d50;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h24f; din <= 32'ha32d3987;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3cc; din <= 32'h8cd66c87;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b0; din <= 32'hb5506e96;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h131; din <= 32'h4ebf7839;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h197; din <= 32'h5270ee15;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c2; din <= 32'h80a6b5b4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h018; din <= 32'h0e2c1fa3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c6; din <= 32'ha7a98043;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h253; din <= 32'hdbec4498;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c5; din <= 32'he804f5e5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2a8; din <= 32'h4cfd85e6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2cb; din <= 32'h722cb078;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h374; din <= 32'h5c81a9ad;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h306; din <= 32'h2ded1cee;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h037; din <= 32'ha8295db0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h238; din <= 32'h6889d421;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h359; din <= 32'h1bdceb49;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h19e; din <= 32'hc7532bc1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h333; din <= 32'h7b6521b7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h004; din <= 32'hdc28db9f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a9; din <= 32'h9d7e88f8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c3; din <= 32'h2942e8ef;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h199; din <= 32'h1c6a4475;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h023; din <= 32'hafb1aa61;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h058; din <= 32'h62e7bb80;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3bd; din <= 32'h6edda060;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h024; din <= 32'hbeb62f98;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3bb; din <= 32'ha1e2c1b9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h17c; din <= 32'h2e4bf5e7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h393; din <= 32'h9bd5eed0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ff; din <= 32'hecdff9c5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h179; din <= 32'h4b05034e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f7; din <= 32'h9904c28f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b7; din <= 32'h505d4230;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08d; din <= 32'h2abc7bb9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e9; din <= 32'hd7c6b576;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c1; din <= 32'h0b0665b2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c4; din <= 32'h7a6e3707;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ec; din <= 32'h10dc9608;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c6; din <= 32'h6aa14a1a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h286; din <= 32'h32722712;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h207; din <= 32'hc5aa586e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h229; din <= 32'h74c7922b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f3; din <= 32'h0f47f304;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d8; din <= 32'h1c325920;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h234; din <= 32'h1855d97a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1fa; din <= 32'ha631fbc8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h384; din <= 32'h4a80c6c3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b7; din <= 32'h6cb43dfb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0da; din <= 32'hde079f54;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h12c; din <= 32'h1ba7f9a7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h377; din <= 32'h43c12856;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h330; din <= 32'h324199dd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h14e; din <= 32'hff26a70e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h232; din <= 32'hde3cc60f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h367; din <= 32'h9e7b1ed0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h117; din <= 32'h19e02ffb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h216; din <= 32'hba27d9a0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h09f; din <= 32'hf06fe077;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d1; din <= 32'h0ea3e44e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h220; din <= 32'h66541038;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h010; din <= 32'h92a754fd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h077; din <= 32'h7df544ab;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h234; din <= 32'h5b017dd2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ef; din <= 32'hea52e9b2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0fc; din <= 32'hd22af72e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h109; din <= 32'h27433e08;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a6; din <= 32'h0ca0c555;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h334; din <= 32'hb06b46db;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h384; din <= 32'heb37c1f2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d0; din <= 32'hce6f09fe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ce; din <= 32'h87434abe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h10c; din <= 32'h24bf68da;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0fa; din <= 32'hf0c9f188;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h225; din <= 32'h71fc15f5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h303; din <= 32'hdb653339;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h246; din <= 32'h25ff502f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ff; din <= 32'h41da7eb3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h334; din <= 32'hfd348b23;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h159; din <= 32'h7b7ba27b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b6; din <= 32'hebf95f25;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ad; din <= 32'hf1490e09;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2af; din <= 32'h7636d28a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h060; din <= 32'hd2b748f6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h182; din <= 32'h3ae0f3ef;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h33d; din <= 32'h9b9acc6c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h01f; din <= 32'h53d85d1a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f3; din <= 32'habf775f2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ab; din <= 32'hccd4aef7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h295; din <= 32'hccb1d1e6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h335; din <= 32'h1b893eb2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e1; din <= 32'h4a351631;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h328; din <= 32'hb3237fbb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h01c; din <= 32'h2654f578;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22c; din <= 32'hf6898d5e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2bb; din <= 32'hb1f0590b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h019; din <= 32'h97012e9d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ce; din <= 32'hea381e3c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h387; din <= 32'h4dfad75e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h046; din <= 32'h2e60dfc3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c1; din <= 32'h05d8fa33;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h280; din <= 32'h28ffe439;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h17b; din <= 32'h9f665286;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ec; din <= 32'h9659f381;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h36a; din <= 32'h8e6a5a8e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h115; din <= 32'h16b8d965;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f6; din <= 32'h33504e98;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37b; din <= 32'h5e569383;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f3; din <= 32'he87ada51;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ae; din <= 32'h5d7f2415;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37e; din <= 32'he02a2324;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h201; din <= 32'hbd6b8fa8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h159; din <= 32'h05708755;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b4; din <= 32'h7e20a8b9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c9; din <= 32'hcb937991;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d1; din <= 32'hedb22404;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e9; din <= 32'h8c47f2ec;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a8; din <= 32'h896fee74;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d8; din <= 32'h89f58e65;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h069; din <= 32'hc1bc1c8b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c3; din <= 32'h434095e3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b5; din <= 32'h3d8fdd70;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d1; din <= 32'ha77f2d37;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h33d; din <= 32'h3e100fec;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h216; din <= 32'h46af0ff4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c2; din <= 32'h4985ec6b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1fa; din <= 32'h70fab136;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3dc; din <= 32'h5cc149b5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h12c; din <= 32'he3a6d6f4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3be; din <= 32'hac2bf194;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1fc; din <= 32'h2637ee0f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16e; din <= 32'hfe6f2e6a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h120; din <= 32'h52ab1547;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2af; din <= 32'h1e6de8e9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d8; din <= 32'hb54fbb29;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2a1; din <= 32'h52792dcc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h19c; din <= 32'hf0578092;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h04c; din <= 32'hd4e41cd5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08b; din <= 32'h1aebccda;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h072; din <= 32'h237567a9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d3; din <= 32'h16aef668;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1eb; din <= 32'h15b2e911;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d7; din <= 32'h562eec91;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h392; din <= 32'h9db3f453;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h29a; din <= 32'hce814d1c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h32b; din <= 32'h0f9d6e16;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ba; din <= 32'h4757780e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h07c; din <= 32'h5dd5f321;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h055; din <= 32'h2c21b128;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23f; din <= 32'hbced0545;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b5; din <= 32'hd9eb8536;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0cf; din <= 32'h35dc1870;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h04b; din <= 32'hce08ca44;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h317; din <= 32'h8d7a1b5b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h083; din <= 32'hda5e8a29;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h008; din <= 32'h729583ff;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h160; din <= 32'h33792436;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h19d; din <= 32'hb49a9776;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b5; din <= 32'hb6870644;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h29d; din <= 32'h39e6a69e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00a; din <= 32'h0d6e8146;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a2; din <= 32'hace987b5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00d; din <= 32'h8bc3736c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h261; din <= 32'hce1b20c7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f1; din <= 32'h7e4c7c2f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h035; din <= 32'ha10e279a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h03c; din <= 32'h2b6fd19a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18f; din <= 32'h3ca02c98;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h367; din <= 32'h9e304c1f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h27f; din <= 32'h14940b95;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b6; din <= 32'h3c1f972d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d8; din <= 32'hf79a1dab;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a3; din <= 32'h389690ad;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h28c; din <= 32'h9884fcc1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0af; din <= 32'h090a0481;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1fa; din <= 32'h67a0f0ea;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3bb; din <= 32'hf390c1e2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d8; din <= 32'hcadda9a6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h253; din <= 32'h92231f92;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16b; din <= 32'h2183153a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h33c; din <= 32'hff275ed6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a0; din <= 32'h12561d13;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h399; din <= 32'he418d77d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h367; din <= 32'h7f40fbd3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h115; din <= 32'h8dbbaec7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22c; din <= 32'he8b73954;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f9; din <= 32'hbb97c9d2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h310; din <= 32'h97b3f185;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h150; din <= 32'hbd89a29c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f6; din <= 32'hdae197da;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h273; din <= 32'h04ce9f82;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ff; din <= 32'h482e7aec;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f7; din <= 32'hcc2e4bfa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ab; din <= 32'hffa0e67d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h367; din <= 32'hf2b9299f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h21c; din <= 32'hf486109a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d0; din <= 32'h5b26479f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2bc; din <= 32'h58c864f3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ef; din <= 32'h7fc11798;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b4; din <= 32'hea6da9cb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37a; din <= 32'h36ff9395;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h36c; din <= 32'h6bf18bfa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c4; din <= 32'h31d107ba;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f1; din <= 32'h16f1a0c3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f4; din <= 32'h5019dbc5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a9; din <= 32'hfb4b5093;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18e; din <= 32'hd8c21d8c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h396; din <= 32'h81a8975a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h34d; din <= 32'hebf7e254;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31e; din <= 32'h14fa69e3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c4; din <= 32'h8e4014d6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h111; din <= 32'h59263c9c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h09c; din <= 32'h949bf477;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h398; din <= 32'hceda03fe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h318; din <= 32'h92a88e1e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h050; din <= 32'h28435e31;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h39f; din <= 32'hef837a98;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3de; din <= 32'h45bef185;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a3; din <= 32'h77374b14;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h184; din <= 32'h0a3afb0d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a1; din <= 32'h0c11cc49;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h163; din <= 32'h2e8064de;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h346; din <= 32'h38b45e21;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h347; din <= 32'hb76ddd48;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h173; din <= 32'h126ec2f8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b5; din <= 32'h1c8db029;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h32f; din <= 32'hb49ecaf5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h102; din <= 32'h6d424029;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h334; din <= 32'h80a3fd45;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h314; din <= 32'h439b18d4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ec; din <= 32'h625fd92f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h316; din <= 32'h3686cd0f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0bd; din <= 32'h2cc3c5fb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h20a; din <= 32'h30e81dae;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d7; din <= 32'h627e4e89;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h221; din <= 32'h42fdc59b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b8; din <= 32'hd1b64e50;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a7; din <= 32'h24e58381;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h27f; din <= 32'h0e9d85f6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f9; din <= 32'haf70b1d8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h15a; din <= 32'h2ad3c13a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ef; din <= 32'h186fa140;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f9; din <= 32'hcafc9463;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h02f; din <= 32'hccfc5c6c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h17a; din <= 32'h9436258b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h131; din <= 32'h54183727;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h219; din <= 32'h57bfd16e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h33b; din <= 32'h53c572e2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c7; din <= 32'hf89fff8e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h268; din <= 32'h30e090c3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h257; din <= 32'h01ee1b46;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ba; din <= 32'h686fd830;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2fa; din <= 32'h195bfcce;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h29a; din <= 32'h98b01b99;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h10f; din <= 32'hebb49673;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h362; din <= 32'hac2e6624;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a0; din <= 32'hd7366ae7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h127; din <= 32'hb725400a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h29f; din <= 32'hbe21c770;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e2; din <= 32'h1245ac5c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h114; din <= 32'h8e691af7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h192; din <= 32'hc0aebc6c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d4; din <= 32'h4ba3ff57;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18a; din <= 32'hbf0801de;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a4; din <= 32'h4499c873;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e2; din <= 32'hb22ee3a6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38c; din <= 32'h2148104d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h079; din <= 32'hb3b453c4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0cf; din <= 32'h110b9f7f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h399; din <= 32'h05263325;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3fe; din <= 32'h92a57aff;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h081; din <= 32'h0844b6f9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d3; din <= 32'h685a7a9b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h084; din <= 32'h8264067c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38e; din <= 32'h90b694f7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h113; din <= 32'h1743902a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e2; din <= 32'h8584293b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ee; din <= 32'h00689192;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00d; din <= 32'h85bfed4d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h016; din <= 32'h25302ac5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0cd; din <= 32'he0bed4d0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b3; din <= 32'hf5c8d6e6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b4; din <= 32'h9f47e76d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h305; din <= 32'heb367558;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h28d; din <= 32'h025569d7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c7; din <= 32'h032a7197;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h297; din <= 32'h021caffe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c5; din <= 32'h5bc757ab;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e5; din <= 32'h83c0d036;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b6; din <= 32'h71f5a10c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h231; din <= 32'h837bfa11;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h125; din <= 32'h18244db9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h15e; din <= 32'h60efa942;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h097; din <= 32'h603ce2a5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e6; din <= 32'h10e4da04;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d2; din <= 32'hfeb808fb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h285; din <= 32'hf5874d0a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2fb; din <= 32'hafa49caa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h09b; din <= 32'ha2af6d2e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h367; din <= 32'hffc15f5b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c0; din <= 32'h44ed177b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h06c; din <= 32'h36739410;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c1; din <= 32'hb01944bd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h323; din <= 32'h845c51ed;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h129; din <= 32'h512ce109;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b2; din <= 32'ha8f16c2a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h245; din <= 32'he20c65d5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h293; din <= 32'h7517b80d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h12c; din <= 32'hc0b8149f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a1; din <= 32'h8b583828;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e8; din <= 32'hdf034c87;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38d; din <= 32'h4b0072a9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h29d; din <= 32'hf82e5b41;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b0; din <= 32'h502d13c7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h352; din <= 32'h0495642f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f0; din <= 32'hc468a143;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h373; din <= 32'h1a0dc2c2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h05a; din <= 32'h932f33ca;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h20b; din <= 32'h0a581df8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h10e; din <= 32'h40bbb011;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h192; din <= 32'h89695958;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08b; din <= 32'hb6205e90;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d6; din <= 32'hfe511745;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h17b; din <= 32'h69e52cfe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37f; din <= 32'hbe0ba911;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h088; din <= 32'h0b7c269a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h351; din <= 32'h8f403ba1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b9; din <= 32'h2d56ea4a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h33f; din <= 32'h3416bba7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h066; din <= 32'hdc37231c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ff; din <= 32'hefa26187;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0af; din <= 32'haa35b073;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h031; din <= 32'h9361464a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h201; din <= 32'h7891069a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h029; din <= 32'h87423eb8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h109; din <= 32'had6d89f2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d1; din <= 32'h6a5f5faa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h356; din <= 32'h72ebe8a5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h322; din <= 32'hf9445dee;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h128; din <= 32'hcbcc93ff;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2da; din <= 32'h991781f9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a9; din <= 32'h35e11dc9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18a; din <= 32'he06bb40c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h042; din <= 32'heb5924dc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h157; din <= 32'h58a4aeea;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h105; din <= 32'h2bedc9a7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h378; din <= 32'h6d9c3991;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h231; din <= 32'h6494eeef;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h224; din <= 32'heaf2e358;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1fa; din <= 32'hd2c8e4eb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h03f; din <= 32'h6599f0ae;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e6; din <= 32'h643d15e9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c6; din <= 32'hab35db3e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h10a; din <= 32'h065d9d34;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h351; din <= 32'h01e84ef1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h006; din <= 32'ha5819f55;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h062; din <= 32'hfeb18c01;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h27e; din <= 32'h975e1947;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37c; din <= 32'h05d3d582;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00b; din <= 32'h66b45dab;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h395; din <= 32'h882cc277;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b0; din <= 32'h4341151a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1bf; din <= 32'h717186bc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h139; din <= 32'h192e5ab6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h389; din <= 32'h8c996a2a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a0; din <= 32'h7828c970;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h351; din <= 32'h0d7c361b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ac; din <= 32'hb578b45f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h058; din <= 32'he027cd4d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d4; din <= 32'h5f4ff6b7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h30c; din <= 32'h47ff09a9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h061; din <= 32'h0a94c0b2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h177; din <= 32'habbc265a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h055; din <= 32'h3af7b8d7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h165; din <= 32'he422aa1e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h02e; din <= 32'h9aa55ca1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d6; din <= 32'hffa8d410;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d0; din <= 32'haceaed9c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h104; din <= 32'ha59c8424;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h116; din <= 32'h21a1b0ae;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0af; din <= 32'h2cbf139b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h016; din <= 32'h100ac447;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h312; din <= 32'hc5a1da68;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h058; din <= 32'he058001f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d6; din <= 32'h5274f255;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0df; din <= 32'h3329cbae;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h372; din <= 32'h7212af50;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h058; din <= 32'ha95576e8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16c; din <= 32'he9a268a6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ab; din <= 32'h613a3abd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a2; din <= 32'h4e9fdf35;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h268; din <= 32'h6f70a801;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0dc; din <= 32'hb6214c76;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a4; din <= 32'he238d762;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h171; din <= 32'h0bcec6b1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c3; din <= 32'h32c7df6c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h12c; din <= 32'he5b3a96a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h30e; din <= 32'h615bee7f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16a; din <= 32'hf509be0c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h015; din <= 32'hf4e9b0b0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h02d; din <= 32'h8ab4399f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c7; din <= 32'h2dfef456;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h227; din <= 32'h9cafe636;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h070; din <= 32'h8cd55f31;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h213; din <= 32'hf19eeccf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h283; din <= 32'h912c65f3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h069; din <= 32'h60b2e3a7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h283; din <= 32'h99d28bf9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16d; din <= 32'h065f0e75;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h141; din <= 32'h2871251a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2eb; din <= 32'h03886424;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b1; din <= 32'h701d208f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08e; din <= 32'h337b5be8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h205; din <= 32'h2f68385b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h046; din <= 32'h9a13933e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ef; din <= 32'h2c7eb56a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h33b; din <= 32'h49da90a6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1df; din <= 32'h673ad5c9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h046; din <= 32'hd645e286;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h093; din <= 32'h5959b225;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ad; din <= 32'h9f99dad0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h39e; din <= 32'h15feb2e6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2a1; din <= 32'he7afe036;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h26d; din <= 32'hce4b1f2f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h370; din <= 32'h1aca5403;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h351; din <= 32'hf26002ee;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c4; din <= 32'hf3254ba7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ce; din <= 32'h699b3736;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h336; din <= 32'haa7f47ba;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ab; din <= 32'hd9d09be3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h229; din <= 32'h1082e92d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h107; din <= 32'ha25b46a4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h19f; din <= 32'h061e299e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f9; din <= 32'hf0c4d24a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h158; din <= 32'h530d920b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ae; din <= 32'h4c677bdb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e7; din <= 32'h58a82c39;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h076; din <= 32'haa21c563;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ba; din <= 32'h6601f400;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h200; din <= 32'h358432cb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2bc; din <= 32'hd0c9ef42;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ae; din <= 32'hfe858c31;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h095; din <= 32'hf3a88dd7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h333; din <= 32'h5c6d26a8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h261; din <= 32'h1ce7bbdd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h219; din <= 32'hacf14bc8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h333; din <= 32'h7854890f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ac; din <= 32'h631b9370;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h01a; din <= 32'h232b5213;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h35f; din <= 32'h55adbcaf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h071; din <= 32'hd85453c0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a6; din <= 32'hd20c086a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e1; din <= 32'h798a2aa1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h260; din <= 32'h08247260;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h03a; din <= 32'h81193810;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3fe; din <= 32'hef8ec073;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31d; din <= 32'hd5181577;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d7; din <= 32'ha663a1bc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h187; din <= 32'h7c50a154;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16c; din <= 32'h3c96088c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h11e; din <= 32'h64026939;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h024; din <= 32'h98d37694;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h28e; din <= 32'h3350ee0e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h093; din <= 32'h77db4692;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0fd; din <= 32'h7e4792f7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e6; din <= 32'h315b85ad;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a6; din <= 32'h4cccfb33;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1cf; din <= 32'hae7c6aff;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e5; din <= 32'h75cf2c6b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ca; din <= 32'h290b8712;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h24a; din <= 32'h7780532d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h264; din <= 32'hd759ad6d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3dc; din <= 32'had2f9440;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d8; din <= 32'h843abe01;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h074; din <= 32'h232876af;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h142; din <= 32'h1bb70605;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e2; din <= 32'h355ef623;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h228; din <= 32'he856d1b0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h239; din <= 32'h36447015;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a0; din <= 32'hcc62af03;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d3; din <= 32'hc348e552;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h25b; din <= 32'h4b1808d8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e3; din <= 32'h0b7878f4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c5; din <= 32'h89860f86;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ad; din <= 32'h6f340a19;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h268; din <= 32'he08af7c3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h392; din <= 32'h496a8871;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h180; din <= 32'hd7dd91a8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h277; din <= 32'hdfd4527e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h13b; din <= 32'heb514f49;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h176; din <= 32'hf869290f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18f; din <= 32'h24ba2dd7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h002; din <= 32'h606c8562;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h14c; din <= 32'heb7537d5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2dc; din <= 32'h446753fe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h217; din <= 32'hd64fdb7f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a0; din <= 32'hc62cdd34;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d7; din <= 32'ha3a89b46;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ab; din <= 32'hf41204ac;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h197; din <= 32'hc3a4118e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2cd; din <= 32'h2fdec321;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h121; din <= 32'h2d87444c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c7; din <= 32'h5c6cd94f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h262; din <= 32'hfb52d744;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37d; din <= 32'h0638ed16;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h20a; din <= 32'ha17cd141;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1cf; din <= 32'h0ad8e518;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23b; din <= 32'hd6bce0ed;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h159; din <= 32'h48d96826;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h143; din <= 32'ha421ce8b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d9; din <= 32'h4f4d2dbd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f0; din <= 32'h22086382;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a9; din <= 32'h94aa6e62;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h03a; din <= 32'hc76d5d34;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0fa; din <= 32'h171da0d9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h30f; din <= 32'hfe86c2e4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h360; din <= 32'h882c54d8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h248; din <= 32'h3795feb4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h282; din <= 32'h17ab4a35;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00e; din <= 32'ha1fb0ac7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h084; din <= 32'h7c6bf113;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h093; din <= 32'h53bf252c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h293; din <= 32'h0ffd403f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h24c; din <= 32'h0ff20371;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c2; din <= 32'h98cabd46;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ed; din <= 32'h4b11bdd6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22a; din <= 32'h954f4d74;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h287; din <= 32'h339a6669;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h14e; din <= 32'h12692036;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h167; din <= 32'h1fdbe3fd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h21e; din <= 32'h5d02face;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h04f; din <= 32'h8a0fd98a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h10f; din <= 32'hbdd9b945;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h108; din <= 32'h77566634;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e0; din <= 32'hd4b7d8e8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h084; din <= 32'h6db59947;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h100; din <= 32'hfd692a9f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h29c; din <= 32'ha6355156;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h316; din <= 32'h1f47b73f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f1; din <= 32'he978e962;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h182; din <= 32'hcb22d639;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h250; din <= 32'hf6244103;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h373; din <= 32'h67ef7a13;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h318; din <= 32'h95527755;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c3; din <= 32'h20ddd064;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23e; din <= 32'h001a5621;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h29c; din <= 32'hccd57e5a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h376; din <= 32'h47bfa6d4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h19b; din <= 32'h0f216bcb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1be; din <= 32'h2b160722;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e8; din <= 32'hb42db15c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23b; din <= 32'he26eb67e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h080; din <= 32'h6b52ff8d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f9; din <= 32'h987daab9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31c; din <= 32'hb57f9edd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h26e; din <= 32'hd7e02980;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a7; din <= 32'h13d694b9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h383; din <= 32'h0709f261;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h39f; din <= 32'h2df6e514;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2a9; din <= 32'hb6a4b840;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h266; din <= 32'h17e8fd57;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d5; din <= 32'h999898c5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23d; din <= 32'h0a991ee8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h051; din <= 32'h843934de;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h335; din <= 32'h41764694;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0da; din <= 32'h090b0637;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f5; din <= 32'h19fb7341;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h15e; din <= 32'hd0e8ee29;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3fb; din <= 32'h1c7472c4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h12b; din <= 32'h56cd5e93;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h02e; din <= 32'h618f9efa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h067; din <= 32'h03bfc437;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h170; din <= 32'hb5833e9e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h333; din <= 32'hf3d69310;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h081; din <= 32'h7ad8903d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h099; din <= 32'h554f0e95;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h339; din <= 32'h6fc9c546;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h003; din <= 32'heb2a6466;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16d; din <= 32'h70cd9a54;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h081; din <= 32'h101a541d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h27b; din <= 32'h3e52f520;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h32f; din <= 32'h9e648ae5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h239; din <= 32'hda7e0437;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h30d; din <= 32'hc2bb1c19;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h17c; din <= 32'hfed54a81;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h357; din <= 32'h505ae374;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h311; din <= 32'h86f5ca26;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b5; din <= 32'h8020ed24;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h30d; din <= 32'h02287f6e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h124; din <= 32'h56f019e1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h227; din <= 32'h73eb44eb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18a; din <= 32'h69e811c8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h203; din <= 32'h0f577b1e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h283; din <= 32'h5513ffea;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b8; din <= 32'hb50c85ad;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f0; din <= 32'h35c6e319;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b9; din <= 32'h1c0b12fa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h253; din <= 32'h366f8067;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h211; din <= 32'h3cce0fb0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h194; din <= 32'h76ba1c99;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h181; din <= 32'hab0d26cf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h271; din <= 32'h47a7df39;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ae; din <= 32'h38173151;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22b; din <= 32'hbf4b444e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c0; din <= 32'h78eef496;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c6; din <= 32'hc5e7e5d6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h022; din <= 32'h8c6975e0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h300; din <= 32'h23c8d0c6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h288; din <= 32'h83830d10;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2a1; din <= 32'h8d2d1643;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h28d; din <= 32'h6f3f2ee2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f0; din <= 32'h99447f4f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h21e; din <= 32'h163180b4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23e; din <= 32'h2ebc47d5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h27e; din <= 32'h142433af;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h15a; din <= 32'h34b02a90;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h20b; din <= 32'h01a45f9e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1cc; din <= 32'h523563c8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h203; din <= 32'h8885ab95;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c4; din <= 32'h7594ac82;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h115; din <= 32'hd73d52d7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a4; din <= 32'h8444b435;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h074; din <= 32'heb449ad2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h353; din <= 32'hdb052fa2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h216; din <= 32'h97c21f73;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h216; din <= 32'hfea25f2a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h01f; din <= 32'h483db685;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f7; din <= 32'h14997081;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e4; din <= 32'h3fbda03f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h157; din <= 32'hbe874ba1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ec; din <= 32'hd0599529;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ee; din <= 32'h724d23f6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38d; din <= 32'h64c82f35;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ab; din <= 32'hb634b7cf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d3; din <= 32'hbcb48b61;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h224; din <= 32'h5407dbc8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d5; din <= 32'hcbe9e18f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h048; din <= 32'h6954048c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h389; din <= 32'hfc300d32;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c9; din <= 32'h62dabc07;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h01e; din <= 32'h0887872b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h231; din <= 32'h02e1bef7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h20d; din <= 32'h522b5a93;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h13d; din <= 32'hfd8b9b64;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h272; din <= 32'h52615401;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h055; din <= 32'ha83d7c82;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h100; din <= 32'h27fc97f9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h19c; din <= 32'h0b2361a1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h14c; din <= 32'he789b252;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f9; din <= 32'h556fa33e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b9; din <= 32'ha18ab8bf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h381; din <= 32'h067a9aca;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h24e; din <= 32'h093ad3e7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1fe; din <= 32'h832f032c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f9; din <= 32'h8e025299;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f4; din <= 32'h74df7b69;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a1; din <= 32'h9777259a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h289; din <= 32'h2435ae96;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a8; din <= 32'hb02788fd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h177; din <= 32'ha954dca4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ce; din <= 32'ha4191b92;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b2; din <= 32'hb360955c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h314; din <= 32'h3434dbd5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e9; din <= 32'ha656b9f0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b1; din <= 32'h3d777fa5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ac; din <= 32'h7ae87ef6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38d; din <= 32'hc130f4fc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h005; din <= 32'h3f1679ab;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h267; din <= 32'hafd25773;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h264; din <= 32'hf56e1781;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h12b; din <= 32'hb4d8583e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2be; din <= 32'h66b08bfe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h32f; din <= 32'h52627642;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h275; din <= 32'ha9a8b471;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h289; din <= 32'h698d72d9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38b; din <= 32'h47afe492;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h387; din <= 32'hcd06fd17;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f8; din <= 32'h64043743;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0bc; din <= 32'hdaf57afa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b8; din <= 32'hbb68cf69;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c8; din <= 32'h64bf79bb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h17d; din <= 32'h23a4ffdf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h359; din <= 32'hd63dc808;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h049; din <= 32'habbeeb19;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h10a; din <= 32'h963cb356;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3fe; din <= 32'h6e662304;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c6; din <= 32'hf5e78d50;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h390; din <= 32'h00ac816b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h230; din <= 32'h91eee5b3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h059; din <= 32'hb4cfab41;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h366; din <= 32'h5f7ac4c9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h111; din <= 32'h2defdefe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ed; din <= 32'h92326aa1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h278; din <= 32'h73380e26;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h15f; din <= 32'h767c472a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h084; din <= 32'hf8615c33;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c2; din <= 32'hde34e75d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h262; din <= 32'h32d69095;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2bb; din <= 32'hd2deb675;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h297; din <= 32'h3ef29e08;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h125; din <= 32'h16a5ada4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0cc; din <= 32'h2cd700e3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ff; din <= 32'h22a2f34d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h172; din <= 32'h7d221d22;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2fa; din <= 32'hb6030221;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ed; din <= 32'hb8f15566;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h318; din <= 32'hed6eac09;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h20d; din <= 32'hdffa81ec;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h092; din <= 32'h6837f33b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h359; din <= 32'h7d52d3c5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h391; din <= 32'he7ebdcb4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h112; din <= 32'h7536b151;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2af; din <= 32'ha0a0db3e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h160; din <= 32'h327fee72;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h29b; din <= 32'h7e5a1c7d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f0; din <= 32'ha2283d80;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h072; din <= 32'h249f60e6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2de; din <= 32'h2c50d85b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31e; din <= 32'hf27d9fe5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h033; din <= 32'hf5c23bc9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b5; din <= 32'hbd4e30d1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31a; din <= 32'h60db3101;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16c; din <= 32'h7ae75106;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h256; din <= 32'hb1ed5fc7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h184; din <= 32'h24fd563c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b2; din <= 32'h7d895a57;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h164; din <= 32'h77d3a908;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h28e; din <= 32'hec33caec;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2da; din <= 32'he6107e57;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h05a; din <= 32'h448e1c00;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h12d; din <= 32'h6609142e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h054; din <= 32'h79049bac;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b5; din <= 32'hff799e36;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22c; din <= 32'h42d59cf7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b7; din <= 32'h7331cf45;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h24d; din <= 32'h7a4c0e78;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f8; din <= 32'h821922ca;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ec; din <= 32'hb178b3af;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h382; din <= 32'h8f1ae5a6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h226; din <= 32'hdab795db;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b0; din <= 32'h3d2b69e5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h342; din <= 32'h2995efba;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a8; din <= 32'h7e1a9204;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h311; din <= 32'hac4b8b0f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h076; din <= 32'h26fff48d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3cd; din <= 32'h7539c0ea;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h07f; din <= 32'hc728dc72;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h212; din <= 32'hdac09a8e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0bd; din <= 32'h978c1f50;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2cc; din <= 32'h70742a4b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h103; din <= 32'h1cfaea84;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h24a; din <= 32'h0c04d6ca;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h30d; din <= 32'h1f7f7be4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ca; din <= 32'h40fd4aaf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h303; din <= 32'hcc382063;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b7; din <= 32'h27ceb9e1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h146; din <= 32'h98fb14c9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h35f; din <= 32'h5581ad20;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h229; din <= 32'h11487879;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2a2; din <= 32'ha4aa9f55;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h389; din <= 32'h3e0f2678;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h32a; din <= 32'hd1071ec2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d1; din <= 32'h0e3a924c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h148; din <= 32'hce015512;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h32b; din <= 32'hfcb005de;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2a7; din <= 32'h3fcd09f7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1cd; din <= 32'hbb907e98;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h314; din <= 32'hf664da16;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h142; din <= 32'h22ac7c99;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h376; din <= 32'hf7673444;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1bd; din <= 32'haafa69f7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h193; din <= 32'h43c8b322;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h169; din <= 32'hb67ccbb2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h197; din <= 32'h00e79ae8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h33d; din <= 32'h1c200cd1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h217; din <= 32'h90dba40d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e5; din <= 32'hda62334b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h191; din <= 32'hbe6ceba8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e5; din <= 32'h328d5a34;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a5; din <= 32'h5f1cccb8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b9; din <= 32'h9755ec40;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h238; din <= 32'h1e475fc8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23d; din <= 32'h58142e38;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d6; din <= 32'hc6c1ffdc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a4; din <= 32'h9a9730b3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h018; din <= 32'h188dd089;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a6; din <= 32'h5afb28fc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h053; din <= 32'h05d7d336;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f3; din <= 32'h53de9737;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h332; din <= 32'hc2827c90;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b0; din <= 32'haa28fb2f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h297; din <= 32'hb3b50bbe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2db; din <= 32'h2f26aa4c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ea; din <= 32'h1e69ba90;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h005; din <= 32'hfaa3b793;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h020; din <= 32'hd7c55636;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h34e; din <= 32'hc4f4662e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f0; din <= 32'hf561b5c8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37b; din <= 32'h17b0030c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h367; din <= 32'h211f4a14;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c0; din <= 32'h1efa697f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h289; din <= 32'hce024999;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d6; din <= 32'hb9be07d0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f3; din <= 32'he7435bcd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e7; din <= 32'h3530c909;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h36c; din <= 32'he515dd8b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h188; din <= 32'h531bcf82;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h019; din <= 32'h0788a3a7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h221; din <= 32'hd5db6a9c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h094; din <= 32'h32844528;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08a; din <= 32'h565077b2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h087; din <= 32'hfdc7de87;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h380; din <= 32'h2078bb1d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ec; din <= 32'hc1404af0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h268; din <= 32'h0303d5c7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h012; din <= 32'h7d053dd0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b2; din <= 32'h479c3f37;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h10d; din <= 32'he53031ae;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h226; din <= 32'he667e751;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ab; din <= 32'hac71931c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h39c; din <= 32'he40bfb21;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h001; din <= 32'ha1f21b18;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h216; din <= 32'h098f6031;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0fa; din <= 32'hc36b5bb8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h29c; din <= 32'hde34324e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d9; din <= 32'hc83c9cb8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d1; din <= 32'hfd1acc45;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h280; din <= 32'h0a990218;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h249; din <= 32'h33705d8b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c3; din <= 32'ha85a09e5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h158; din <= 32'h447050ad;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c5; din <= 32'h4abe266c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h11b; din <= 32'hd44783c3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h13d; din <= 32'h10652959;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h027; din <= 32'he6454a25;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e0; din <= 32'h4eeb0262;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h35e; din <= 32'h48b1b1d6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h162; din <= 32'he98e33c8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f7; din <= 32'h9503bb52;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37d; din <= 32'he18a085c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b5; din <= 32'hab6e6712;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a7; din <= 32'h06a0f9ff;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h124; din <= 32'h4c770443;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h24f; din <= 32'hdea3e60d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b1; din <= 32'hfdd8cc8e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h388; din <= 32'hb10248e0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e6; din <= 32'hb3a12b6a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c6; din <= 32'h632b6d46;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h04e; din <= 32'h170769b0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h086; din <= 32'hece49982;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2aa; din <= 32'h1f7a962a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h223; din <= 32'h61bf5bd9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e0; din <= 32'h5db146d1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h266; din <= 32'h315fde94;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1df; din <= 32'h62262eec;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h233; din <= 32'hdbf02308;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h181; din <= 32'h56653198;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h04b; din <= 32'h95a12cf4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f3; din <= 32'h30bbdc0f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h178; din <= 32'h7d5ec925;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18c; din <= 32'he967f7f2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16e; din <= 32'ha62b9d77;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37f; din <= 32'hfe8aa4e5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3bf; din <= 32'h98b0eac8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22c; din <= 32'h1d332aa3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h14d; din <= 32'hd80ee405;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00a; din <= 32'ha6dbd47a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h314; din <= 32'hacd7ad67;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1fe; din <= 32'h1794db99;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h10c; din <= 32'hd7c89702;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c3; din <= 32'h53fba1c7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h067; din <= 32'h50b7fa8c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ce; din <= 32'h0b269f41;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h17d; din <= 32'h9378e264;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0fc; din <= 32'h81526187;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e2; din <= 32'h10e2c62c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2fd; din <= 32'h6d17d438;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f0; din <= 32'h5c1c41c5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h24a; din <= 32'h4ff1eb26;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h26b; din <= 32'h46a1216e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h042; din <= 32'h5b735e4c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e5; din <= 32'h52b394e9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0cc; din <= 32'h07c18b10;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e7; din <= 32'h74f56329;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2fd; din <= 32'h9d12e743;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f9; din <= 32'h16deac25;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h160; din <= 32'h42f2c695;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h20f; din <= 32'hb1898d96;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h325; din <= 32'h8497b213;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h276; din <= 32'heb7a008e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c0; din <= 32'h5ea21390;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h385; din <= 32'h212f747a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h137; din <= 32'h98b8b796;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00d; din <= 32'h82616d7f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h170; din <= 32'h63b3ae3b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ff; din <= 32'h8e1003cb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2cc; din <= 32'hf436e8ad;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h339; din <= 32'he1eadeba;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h204; din <= 32'h83c92284;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f4; din <= 32'hfa938731;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00c; din <= 32'hbc397351;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h394; din <= 32'h5d26f9cc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h152; din <= 32'hfbc6ba3b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ed; din <= 32'hd59afbd5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3fe; din <= 32'habad5d82;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h152; din <= 32'h073b8c33;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h13b; din <= 32'h8e1facdd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a0; din <= 32'h52b18c0e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h386; din <= 32'h240a8e5d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h253; din <= 32'hfb55c670;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h315; din <= 32'hbc59c338;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h191; din <= 32'h9896b8e1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h363; din <= 32'h63183644;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31e; din <= 32'h74d2788a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c3; din <= 32'hca5ced34;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e5; din <= 32'h8d688717;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b5; din <= 32'hdce66d6c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b9; din <= 32'hc3b7db8f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h055; din <= 32'h1372b558;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h359; din <= 32'h8095370e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f5; din <= 32'h4c50ccc9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h217; din <= 32'h3b5b59a6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h015; din <= 32'hf5949149;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1cd; din <= 32'h94e7d245;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ba; din <= 32'h36dfcef2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h175; din <= 32'h7328f9e4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h083; din <= 32'hf752a7f6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h054; din <= 32'h0717dd4b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ad; din <= 32'h4b787aa4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a4; din <= 32'h15014af8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f2; din <= 32'hfaadc731;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h002; din <= 32'h176ad833;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h36c; din <= 32'he6ec83db;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h349; din <= 32'he95b9b34;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c8; din <= 32'h7f011c94;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h017; din <= 32'h1f191c97;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h34e; din <= 32'h631ab273;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h06f; din <= 32'hc9010115;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d8; din <= 32'hf6c20454;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ec; din <= 32'h1281749c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h378; din <= 32'h695514a8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18b; din <= 32'ha9f50ee9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a5; din <= 32'h4741ef23;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h390; din <= 32'h01787ce8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h17e; din <= 32'hf7b20155;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h366; din <= 32'hf38e0dbf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h352; din <= 32'h807a4d00;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h32e; din <= 32'h300d9caf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h102; din <= 32'he68af1b9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h022; din <= 32'h0967dc3e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b9; din <= 32'h1ffab26a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0aa; din <= 32'h5ec7c72a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h276; din <= 32'h0cd3c81e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2be; din <= 32'h9b6018eb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ba; din <= 32'hf895d581;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h14a; din <= 32'he898ad4b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b9; din <= 32'habb7a460;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h396; din <= 32'hc4bc53f4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h088; din <= 32'h7999b3fb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c4; din <= 32'h5b0e8668;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h077; din <= 32'h0883af1c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23b; din <= 32'hc2b11c86;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h02f; din <= 32'h26718aff;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c8; din <= 32'he0d08e6b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h365; din <= 32'hecf32e3e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h327; din <= 32'hd7d39e26;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h10c; din <= 32'he9bf0db9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ec; din <= 32'hbe96d1d5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f8; din <= 32'hdf6bce33;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d4; din <= 32'h93ee6286;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h06c; din <= 32'h01de1d8a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3dd; din <= 32'h54bccd9c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h132; din <= 32'h2da71a44;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h240; din <= 32'haeee4175;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h054; din <= 32'hb61cc847;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h009; din <= 32'hf6e4e36c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1dd; din <= 32'h49e4113d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c4; din <= 32'h73fa8a64;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d4; din <= 32'h3b4539ce;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h203; din <= 32'h4f305374;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h278; din <= 32'heb134441;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23b; din <= 32'ha9741c0f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h175; din <= 32'h6f8fac6d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h230; din <= 32'he0ea7ac0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h268; din <= 32'hb8f70a22;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e5; din <= 32'h30e25d93;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f5; din <= 32'h029f5d51;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c2; din <= 32'h3ea02d5e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0fd; din <= 32'hddf5ff04;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h15d; din <= 32'haa80afc1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h219; din <= 32'h05ac4a99;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h145; din <= 32'h6ea3f01d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1dc; din <= 32'he619d2d2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h358; din <= 32'h9775f2ff;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ec; din <= 32'hed74cd8b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h14a; din <= 32'h2d4a0f51;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ca; din <= 32'h7592528e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h34e; din <= 32'h2e6e679b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0be; din <= 32'heeff6a04;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h26d; din <= 32'hc9a76ead;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h394; din <= 32'h486cb9b2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2da; din <= 32'h26b8dee8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c1; din <= 32'hb11d2be6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h25e; din <= 32'hb8ed4c5a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h279; din <= 32'h173d2af4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h191; din <= 32'hc677bd82;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h06c; din <= 32'h06223d1a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h063; din <= 32'hef216158;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h075; din <= 32'hacb66c34;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0bb; din <= 32'h9611a800;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ac; din <= 32'heec7a214;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38d; din <= 32'hc3da5ccb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h27e; din <= 32'h467dbe97;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ba; din <= 32'he7c67c98;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h008; din <= 32'h8eea2c23;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h267; din <= 32'h36950f83;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d7; din <= 32'ha4028875;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h223; din <= 32'h7437e788;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h053; din <= 32'h592aad3c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h146; din <= 32'hd9211489;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b7; din <= 32'h15533e13;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2a5; din <= 32'hbd73760b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h021; din <= 32'h9f8ffbf7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ad; din <= 32'hf0c9bd81;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h246; din <= 32'h5b787c36;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h127; din <= 32'hc58464c4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h06d; din <= 32'had4c2ab1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h035; din <= 32'h140a1b6d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23c; din <= 32'hc6624bd9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h15b; din <= 32'he383e15b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e6; din <= 32'hc1b0fdf5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h058; din <= 32'hb1ad7a20;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b7; din <= 32'h202acedf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2bb; din <= 32'hc535f11a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h251; din <= 32'hfb68e4e8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h15e; din <= 32'he01c1217;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2cf; din <= 32'hab4b8ebe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b8; din <= 32'hed6087a9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ed; din <= 32'hadd9a299;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h25a; din <= 32'hd0a29820;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c1; din <= 32'h152dd4e7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18c; din <= 32'hb70e1acf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h319; din <= 32'ha3bc7090;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h234; din <= 32'h74dd50dc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h088; din <= 32'hb5cdc92c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h143; din <= 32'he4b8c92e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38e; din <= 32'hdec0b03f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h098; din <= 32'hf63f766a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c2; din <= 32'h0762ccf9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e6; din <= 32'h3ce809a9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a1; din <= 32'h8910113b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e1; din <= 32'h755df55f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31d; din <= 32'h1e3bd6d1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ba; din <= 32'h027a817d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h07e; din <= 32'hf487f7a5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h180; din <= 32'h73537011;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h10b; din <= 32'h08518ae5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h086; din <= 32'hb970d79b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a5; din <= 32'h91d6de76;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1cb; din <= 32'hb5686a22;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h152; din <= 32'h0e556db5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h092; din <= 32'h50185fec;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1da; din <= 32'h56ccb65d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b9; din <= 32'h54857e14;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h220; din <= 32'hbef9b085;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d0; din <= 32'h87bd3131;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h181; din <= 32'hf31426a2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h35f; din <= 32'h677ec7e8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c7; din <= 32'hc0e5f742;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3cd; din <= 32'h03c213ee;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38e; din <= 32'hb83fbee6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e9; din <= 32'hac026f47;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h171; din <= 32'h84e39ff1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d9; din <= 32'hb3bc9c84;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c2; din <= 32'hfc047c34;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h04e; din <= 32'h871f7c95;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1de; din <= 32'h83575b49;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e5; din <= 32'h6c0908a2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h02d; din <= 32'h2e27f7f4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h352; din <= 32'h1351bfc8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h264; din <= 32'h5e3b6244;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h21e; din <= 32'h296d3719;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h15f; din <= 32'h0630cbab;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b9; din <= 32'h612bd5c9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h27c; din <= 32'hb300010f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h20c; din <= 32'hb03df8be;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h219; din <= 32'ha3e04190;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2fe; din <= 32'h53b81660;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d7; din <= 32'h272e4c5a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h117; din <= 32'hdf5f6725;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h305; din <= 32'h3a8c89d8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h142; din <= 32'h59341ba7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h25d; din <= 32'h25e121f8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h056; din <= 32'h13bc7ba1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23c; din <= 32'h765ce717;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h287; din <= 32'h64312c34;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h362; din <= 32'h6886b2f8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h066; din <= 32'hf8fa24ae;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h058; din <= 32'hd5778bac;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18d; din <= 32'h15cb7ef8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b3; din <= 32'h73dc6346;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23b; din <= 32'h83f9bc0b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3da; din <= 32'hcdfc53c9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f6; din <= 32'hade283e7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2cb; din <= 32'h3749efe1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h262; din <= 32'h7ec85b24;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h151; din <= 32'h425fdde5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h118; din <= 32'h62dc8732;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h147; din <= 32'h79a7a473;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1de; din <= 32'h28d14b63;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ed; din <= 32'h2a421f16;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f4; din <= 32'h81c0f10c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3cc; din <= 32'h75212b77;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h02e; din <= 32'hcfcc6d83;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d4; din <= 32'h79544d71;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0bd; din <= 32'h768f4bb2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d8; din <= 32'h40ff6193;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h005; din <= 32'ha8420189;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3eb; din <= 32'h76c7e542;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0bf; din <= 32'haf351710;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c6; din <= 32'h165a736b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h15a; din <= 32'h007b1f57;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1af; din <= 32'h340ddf5b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h138; din <= 32'h50924683;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h296; din <= 32'he9623fc5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h03e; din <= 32'h35da2734;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3aa; din <= 32'h5de7f554;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b3; din <= 32'hc38062f6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h255; din <= 32'h0a23e979;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h39a; din <= 32'hf484719f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c3; din <= 32'h8271a684;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a6; din <= 32'h9e5ca726;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ec; din <= 32'he1ac0f40;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d8; din <= 32'hdff28815;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h138; din <= 32'h0023e984;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2dd; din <= 32'h11e8fc0e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h28a; din <= 32'h0550b288;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h340; din <= 32'hf9ef56f0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2fe; din <= 32'h6561752a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h348; din <= 32'he55c1073;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h35d; din <= 32'h079920ae;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h068; din <= 32'h0821aad7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h04c; din <= 32'h27df9601;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d5; din <= 32'h061bcd61;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h06d; din <= 32'h4a5e650d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0dc; din <= 32'hd96d6f56;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3dd; din <= 32'h18340333;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h09c; din <= 32'h745035ce;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e8; din <= 32'h349a4e1a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h399; din <= 32'h020a3abc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b2; din <= 32'hfb67be82;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0bf; din <= 32'h80c5a4a5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h153; din <= 32'h6377e7b6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h310; din <= 32'h24c84a6e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h160; din <= 32'h41607477;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h12b; din <= 32'h63f929c8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c6; din <= 32'h29c6245c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c7; din <= 32'he909c177;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e2; din <= 32'h352c4159;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b6; din <= 32'h637a1bc0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h248; din <= 32'hf2a4e639;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b5; din <= 32'hdca89229;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0fe; din <= 32'h21e360d7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h316; din <= 32'h9d9a0151;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h33e; din <= 32'hb6862e0c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e7; din <= 32'h54da60aa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e1; din <= 32'h0e522986;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1bd; din <= 32'h12b3a86e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h04d; din <= 32'hc5ec15fb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h393; din <= 32'h5c4c9b03;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h382; din <= 32'he43bcc47;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h160; din <= 32'h5279cb58;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d1; din <= 32'hce69c436;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2a4; din <= 32'hd6e1dc16;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h346; din <= 32'hf5311648;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3cb; din <= 32'h07df76ba;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h146; din <= 32'h0fd4ff65;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f5; din <= 32'h4b946ac2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h383; din <= 32'h7f79bc7d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ae; din <= 32'hb98af2e9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a1; din <= 32'h5936c833;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c2; din <= 32'h7e9196fe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1fa; din <= 32'h9991e86f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h088; din <= 32'h7fd47fb8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h013; din <= 32'h7a8a493c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2a0; din <= 32'hdec43f76;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h156; din <= 32'hd5f76db8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h361; din <= 32'hfd1aedf4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d2; din <= 32'h9a54457e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h369; din <= 32'h81a80cce;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h319; din <= 32'hb211d6c0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d2; din <= 32'ha3deadfd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h017; din <= 32'ha3c73c94;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h164; din <= 32'h0aa003bd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1bf; din <= 32'hbea3fab0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h237; din <= 32'hbaac91f2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h36d; din <= 32'hcfc62256;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h11b; din <= 32'h3c470961;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h189; din <= 32'h472664a0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0aa; din <= 32'hf3a49380;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h200; din <= 32'hc530550d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f3; din <= 32'hf7e662f6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h368; din <= 32'h9cccc465;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a5; din <= 32'hb91b407e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h090; din <= 32'h78aed81a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ac; din <= 32'h8c5f0f81;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h093; din <= 32'h892a7bc0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h344; din <= 32'h9707258b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16b; din <= 32'h29cd0135;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h15b; din <= 32'h439d7f85;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e6; din <= 32'ha2d13611;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f9; din <= 32'h23326df7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f9; din <= 32'h24e76d8b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f7; din <= 32'hf1dd353b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31f; din <= 32'h6b8594e5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h21d; din <= 32'h11bcb107;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2db; din <= 32'hf28ccaa1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h39a; din <= 32'h7f5fe2db;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h389; din <= 32'h0db42deb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b3; din <= 32'h4acb0eb7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h288; din <= 32'hef998cca;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0db; din <= 32'h87bef53f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h366; din <= 32'h0b9e1b15;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h062; din <= 32'h96abf25a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ed; din <= 32'hddc692b2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23d; din <= 32'h2755840e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e6; din <= 32'h831f43f5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h322; din <= 32'h8c5c9f8e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h337; din <= 32'h4acfb4ed;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h19b; din <= 32'h147927cf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37c; din <= 32'h648c3823;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h330; din <= 32'h81218afe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b3; din <= 32'hd846f22a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h260; din <= 32'h7e94212c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c8; din <= 32'h49cf0a4d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h276; din <= 32'hff07b149;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b8; din <= 32'h687ccedc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h343; din <= 32'h8d8db8cb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h089; din <= 32'hc80557c2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h195; din <= 32'h7d6f40ae;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c0; din <= 32'ha04d3067;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c8; din <= 32'h82a34409;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ae; din <= 32'hf4c75137;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c7; din <= 32'hae171e40;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h016; din <= 32'h0700e9dc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h011; din <= 32'haf02286b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h291; din <= 32'ha39ef671;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h375; din <= 32'h937cc8d2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h258; din <= 32'hf30b297d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2bd; din <= 32'hd3fbd476;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b1; din <= 32'hf06c146c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h039; din <= 32'h4bc3acc8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h20a; din <= 32'h2442b1c8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h212; din <= 32'h2012a039;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ac; din <= 32'h01e4cf62;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d1; din <= 32'hcbd5db5b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h21f; din <= 32'h95002bff;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c5; din <= 32'h6e8ecc4c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a2; din <= 32'h533b232a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h161; din <= 32'he5397da7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0db; din <= 32'h94d8e2a8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0eb; din <= 32'h4c99df6a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h03e; din <= 32'hb50010a1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e5; din <= 32'ha256971c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00f; din <= 32'h41801beb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f3; din <= 32'h7bdeb635;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e1; din <= 32'h49c19a1a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31d; din <= 32'h1880dd48;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h325; din <= 32'he39965dd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h382; din <= 32'h6724ba0a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h36c; din <= 32'hfc8e3656;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h14f; din <= 32'hf0b596f4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h338; din <= 32'h00db6883;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h197; din <= 32'hb65d74a7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e6; din <= 32'haf600e8d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ac; din <= 32'hbc0ac611;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h279; din <= 32'h02563207;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h132; din <= 32'hb99b77c3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f8; din <= 32'hc9851f70;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a0; din <= 32'h4eac057d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h060; din <= 32'h7052484a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h271; din <= 32'h56d87fff;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h20f; din <= 32'h46336b61;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08d; din <= 32'h5d51c298;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ec; din <= 32'h4c5cd1de;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d1; din <= 32'h01f69e6a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d2; din <= 32'hcddae9ed;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b4; din <= 32'hfee75779;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e3; din <= 32'h507e5547;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h116; din <= 32'ha276ad68;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h10a; din <= 32'h66026d15;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h11d; din <= 32'h1aa9b04c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d1; din <= 32'hf52819b7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e6; din <= 32'h8818a173;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h310; din <= 32'habbb9247;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08b; din <= 32'h4c417779;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h27e; din <= 32'h5222721b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h303; din <= 32'hb4f59319;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h36c; din <= 32'he0e5b168;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e2; din <= 32'h3e9fd381;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h243; din <= 32'hee742cdd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f3; din <= 32'ha9f71d8d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e5; din <= 32'h3412d1b9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23b; din <= 32'he48c83f7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h21c; din <= 32'hd6195cd1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h02f; din <= 32'hca2395c5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ed; din <= 32'h4affe841;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h003; din <= 32'h1c5b1bc5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h333; din <= 32'h04b96d5c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h087; din <= 32'hdba61830;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h03c; din <= 32'h9636c393;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ba; din <= 32'h89448db5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h386; din <= 32'h6e8c38f6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h046; din <= 32'hf9c4eada;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h388; din <= 32'h42ef2bf7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h380; din <= 32'h9673568e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h12b; din <= 32'h8205ac21;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b7; din <= 32'ha9b67460;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b5; din <= 32'h4789915d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h191; din <= 32'h197136c3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1fd; din <= 32'hb4e96b54;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h15c; din <= 32'h1457c896;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h140; din <= 32'hbc230557;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f6; din <= 32'h6b4eec4b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h360; din <= 32'hb0c5b3e9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h30a; din <= 32'h56b42c45;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h388; din <= 32'h7c760621;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h126; din <= 32'ha5626f0d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h388; din <= 32'h7f2f3ec0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h06c; din <= 32'h35170b61;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ee; din <= 32'h33a20d06;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h158; din <= 32'hb7776eb5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18c; din <= 32'hbccb0e35;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16e; din <= 32'h59e08dad;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16b; din <= 32'he15b2381;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h359; din <= 32'hd77676bf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h12f; din <= 32'h45c0c503;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b7; din <= 32'h69ecadb9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h01b; din <= 32'hff82a74f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h091; din <= 32'h209b3889;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1fb; din <= 32'h485f3638;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0bc; din <= 32'h15f5e794;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d9; din <= 32'h7d6303fc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h26f; din <= 32'h227bd685;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ee; din <= 32'hd815662f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h107; din <= 32'h0da124e2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h394; din <= 32'hf2b9f7f9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ee; din <= 32'he9e6313f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h344; din <= 32'h29799908;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37e; din <= 32'h11aceda8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f3; din <= 32'h0d5ef27e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h353; din <= 32'h4816ad09;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h32c; din <= 32'h15e5a17c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h307; din <= 32'hcda7b04f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ae; din <= 32'h13009b98;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h163; din <= 32'h66d3ec88;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h278; din <= 32'hd25e628a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h235; din <= 32'h318b0a9f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b3; din <= 32'h6bd3e8c3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h127; din <= 32'h54190836;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38a; din <= 32'hd863e6dc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f8; din <= 32'h55ce87e3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c3; din <= 32'hd629f8bb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ae; din <= 32'h0dfcff07;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h03e; din <= 32'hbefe973c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h27a; din <= 32'h88f24eb4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31c; din <= 32'h3a69945b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h017; din <= 32'h6f9e53e1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h325; din <= 32'h5141df7f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h032; din <= 32'ha9971e3d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ca; din <= 32'h9375443d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2cb; din <= 32'hcecb891a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a6; din <= 32'h77b09bd5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h055; din <= 32'h97c21b8f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h095; din <= 32'h11a735b3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e4; din <= 32'h74a3b790;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h01d; din <= 32'h4d3eb836;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c8; din <= 32'h5c5e8392;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h399; din <= 32'hf7330160;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0bf; din <= 32'h07e17a3d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h352; din <= 32'h8cfa6aa5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3da; din <= 32'hab09f7dd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0eb; din <= 32'hf66f07a0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h19e; din <= 32'h281888eb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e9; din <= 32'h59cb24bf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h122; din <= 32'h4140a264;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h310; din <= 32'h982466f9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e2; din <= 32'hafa012cc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h276; din <= 32'h35b32a59;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h026; din <= 32'h455e9094;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ae; din <= 32'h00a3c5ed;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h04e; din <= 32'hc4e4323f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ce; din <= 32'h9a04c8fe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00a; din <= 32'h3d387211;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16a; din <= 32'h3147d43b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h063; din <= 32'h60db545f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c3; din <= 32'hb241a649;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f0; din <= 32'h84d661f9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h147; din <= 32'h1ebcad88;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h30f; din <= 32'h7db6348f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h33a; din <= 32'hb605b4f5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h28e; din <= 32'hc5d386c9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h21a; din <= 32'hd463b22c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d0; din <= 32'hd42e44ff;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a6; din <= 32'h348c7fc6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b8; din <= 32'he87aa8c9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b3; din <= 32'h76c02360;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h369; din <= 32'h2e1f0de4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h254; din <= 32'he6fbb2e6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0aa; din <= 32'hf014aacc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c3; din <= 32'h70bb30c4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c8; din <= 32'h66fbc358;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h21a; din <= 32'h215deb05;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h25d; din <= 32'h482a6177;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08a; din <= 32'h2568bece;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ed; din <= 32'hd5c4e8b8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h267; din <= 32'ha071413f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h284; din <= 32'habf8c233;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22d; din <= 32'ha2dad65a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31e; din <= 32'hc961cbff;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h343; din <= 32'h6971a634;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b0; din <= 32'hbd7ba73b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h014; din <= 32'h8bec3523;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h155; din <= 32'h5a24f1eb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c5; din <= 32'h08f17c69;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h09d; din <= 32'h6ab8ef1e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h172; din <= 32'hfd8d727b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ea; din <= 32'hc8825555;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h277; din <= 32'h9702f64a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h213; din <= 32'h5799b6e8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h363; din <= 32'hd3b54a84;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h15b; din <= 32'he6db12cb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2bf; din <= 32'h527c101e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2cb; din <= 32'h9d168abb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h087; din <= 32'h61e6aa70;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2bb; din <= 32'h26e9f062;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h124; din <= 32'h0820d41c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f4; din <= 32'h02476481;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h36c; din <= 32'h43574d34;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31a; din <= 32'hebd9ede2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h375; din <= 32'ha411fb2c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31b; din <= 32'hec69fc71;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h33f; din <= 32'h5487d35a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h057; din <= 32'hffdc12fd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h168; din <= 32'h249c0a52;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h316; din <= 32'h56a5089d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h112; din <= 32'hb9b4d040;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3bc; din <= 32'h585bb6fd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f1; din <= 32'h773c834a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ac; din <= 32'h7971bb7a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h137; din <= 32'h271634ec;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h33a; din <= 32'h67dbb62e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2cb; din <= 32'hd3fe69d6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2cf; din <= 32'hb0d60a8c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h09e; din <= 32'h14f91e13;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ad; din <= 32'heb23ae6b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h238; din <= 32'h9d859545;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h188; din <= 32'hd350dc0a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ab; din <= 32'h584303d8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h06d; din <= 32'h702ecb07;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22d; din <= 32'ha7583fc3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ca; din <= 32'h29334c8e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37f; din <= 32'ha4a22451;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h351; din <= 32'h147fee00;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h302; din <= 32'h702e4b2a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h040; din <= 32'ha4bf505d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38c; din <= 32'h4ed0a2e5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ce; din <= 32'h8cb7fe08;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h221; din <= 32'h50508ada;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2fc; din <= 32'hde9b2e1f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h03f; din <= 32'h66b48681;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h273; din <= 32'hf831edc4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h07e; din <= 32'h530dfdc3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h13d; din <= 32'he8fff59c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h131; din <= 32'hf291a8bc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h28a; din <= 32'h36fec016;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h11e; din <= 32'h01fc64af;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00e; din <= 32'ha2fd7dd4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h06d; din <= 32'h2162ff23;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18f; din <= 32'h7301b1a0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h113; din <= 32'h6b768c62;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c2; din <= 32'h079c2149;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1bb; din <= 32'hb62bcb87;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b2; din <= 32'he445acdc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ed; din <= 32'h192d48d4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h04a; din <= 32'h2555f9f5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h12e; din <= 32'h9b7d5e9d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h193; din <= 32'h17cd3aa5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00f; din <= 32'h63ed2be9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h312; din <= 32'h13fe49af;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h103; din <= 32'h70d09c4b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h17a; din <= 32'h2ed6e05d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c1; din <= 32'he27ee1cb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2dc; din <= 32'h7b152f12;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1fe; din <= 32'hd3ed8f6b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37b; din <= 32'he01c4e5a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h10b; din <= 32'h7e6789ce;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1aa; din <= 32'hc137bec7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08b; din <= 32'h0c26591b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h160; din <= 32'h269418d4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h15e; din <= 32'hb3783e32;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h20f; din <= 32'h6c508ef6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h314; din <= 32'ha069f255;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a8; din <= 32'hdfb616ea;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h097; din <= 32'hcf2dfd4a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h073; din <= 32'h06d59fc1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38e; din <= 32'h8b77f118;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e9; din <= 32'haa7faadd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h33f; din <= 32'hfdfabe63;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h15a; din <= 32'h2aac1451;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h286; din <= 32'h8f349860;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2df; din <= 32'h7af233b9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h30a; din <= 32'h12f2d792;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h26d; din <= 32'he193adc4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h333; din <= 32'h4acba830;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h373; din <= 32'hc2755c09;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ca; din <= 32'h883db645;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h312; din <= 32'hcafb1718;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c3; din <= 32'h7ca70e62;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h27b; din <= 32'hd80decdd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h105; din <= 32'hb8a80a35;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h140; din <= 32'h8a891491;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ba; din <= 32'h8e67b01c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h313; din <= 32'hb0a2c042;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h234; din <= 32'hd09efffd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e6; din <= 32'h55359ddb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h05d; din <= 32'hcbe30867;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c4; din <= 32'hc4337ceb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h163; din <= 32'hfb46b651;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3bb; din <= 32'hb8bf5ccf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h187; din <= 32'h157db4b6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h052; din <= 32'h6b7f6375;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23d; din <= 32'h803dff83;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h176; din <= 32'h5f53f135;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2de; din <= 32'heaf5bb07;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b1; din <= 32'h27be8b6f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e5; din <= 32'h93663c1d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h35a; din <= 32'hdc5a4758;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c3; din <= 32'ha40d3c37;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h101; din <= 32'h813255c7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h14f; din <= 32'h6172dc8f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h281; din <= 32'h1756a00d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c8; din <= 32'h278704ab;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h269; din <= 32'he968c8b7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2cf; din <= 32'h1d20cb56;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h06d; din <= 32'h14f41811;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h39f; din <= 32'hab417ace;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ec; din <= 32'h0fd660c7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08a; din <= 32'h216bbc7c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h02c; din <= 32'hd1560021;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h123; din <= 32'hc377e73d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h28f; din <= 32'h8c249e3c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h27f; din <= 32'h55eb75b6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h201; din <= 32'h767e11ec;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h07e; din <= 32'h975587b0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3af; din <= 32'hd20e5e49;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e9; din <= 32'h6fcafd90;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18a; din <= 32'h4eb5fcde;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h017; din <= 32'h7320e93a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ce; din <= 32'h9ab9327d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h364; din <= 32'h676f4658;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h288; din <= 32'hb85248f5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h15e; din <= 32'hc538161e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d4; din <= 32'hd84055c2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b8; din <= 32'h3dc41399;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c9; din <= 32'h559bd4e2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ca; din <= 32'hae6fa461;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h07a; din <= 32'h2dea1dbc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23c; din <= 32'hc71c34fe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d6; din <= 32'hc2462b0d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h265; din <= 32'h6289852c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h095; din <= 32'haf3afdde;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f6; din <= 32'h18aabbdc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h166; din <= 32'h5d6554a0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1bb; din <= 32'h33a6d605;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1bd; din <= 32'h9e9f4c8b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e2; din <= 32'h63a7ab69;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h073; din <= 32'h14b3ba06;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a1; din <= 32'hf8296d25;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h129; din <= 32'h7a3afe91;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d3; din <= 32'heddd25d9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c7; din <= 32'h7bb0683c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0da; din <= 32'h6b1a901c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ba; din <= 32'h09a7766d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c4; din <= 32'h78386ff7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h12a; din <= 32'hfaa4b064;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h302; din <= 32'hc399ed64;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22a; din <= 32'h2b0a899b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23b; din <= 32'h15a73fea;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h32a; din <= 32'h1300baac;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h33e; din <= 32'h1679ce4f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h232; din <= 32'ha9c8a860;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3cc; din <= 32'h9f32680b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h030; din <= 32'ha6c6c78d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h028; din <= 32'he3242216;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h076; din <= 32'h381f2e6d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h15d; din <= 32'h258a91bc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e4; din <= 32'h92f72597;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h14b; din <= 32'h3b8c606e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h321; din <= 32'h559676be;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b2; din <= 32'he620781c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h28e; din <= 32'h5be1c99e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1eb; din <= 32'h2370bad5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c5; din <= 32'hd28e9109;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h12a; din <= 32'he0a7a0cf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h269; din <= 32'hd7bbf65f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h27e; din <= 32'h04320ec7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h152; din <= 32'h82ecbab9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d0; din <= 32'h099e7857;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h018; din <= 32'he3b3ccbf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h09a; din <= 32'h9ac05f53;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h259; din <= 32'h9119cf35;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h21f; din <= 32'ha9a049d1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h36a; din <= 32'h6a8c16cd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b1; din <= 32'hef791f74;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h178; din <= 32'h210700cc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22a; din <= 32'h713e8437;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h093; din <= 32'h17b47e36;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h09a; din <= 32'h0c305309;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a8; din <= 32'h3ba93b13;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d2; din <= 32'h97165cbe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h384; din <= 32'h7034995a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ef; din <= 32'hc40e9bca;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h229; din <= 32'h6a6663d9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h274; din <= 32'hbdba6029;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h203; din <= 32'h51983650;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d1; din <= 32'he76445a2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c7; din <= 32'h735adce8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h008; din <= 32'h309b22ff;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f2; din <= 32'h51091dfc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h055; din <= 32'h136b354a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h189; din <= 32'h91b178e4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h296; din <= 32'h1d4f6b3d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ab; din <= 32'hafdcc67f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h25a; din <= 32'h1f8a95a3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h336; din <= 32'h0c3b5383;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h387; din <= 32'h6dc74e27;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h076; din <= 32'h3c103b20;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f1; din <= 32'hf0fb6589;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2cf; din <= 32'h2aabb828;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h136; din <= 32'h81295e5c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f6; din <= 32'hee51e2bb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e2; din <= 32'h40bf65c3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d3; din <= 32'h4a402730;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h28b; din <= 32'hd29ab6d0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e3; din <= 32'h9b6069dd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b1; din <= 32'hd5d427a9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b8; din <= 32'h99f28382;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h06b; din <= 32'h88a25e0f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c4; din <= 32'hf914d1dc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h028; din <= 32'h9c5da801;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ea; din <= 32'h11953f84;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h227; din <= 32'h2d86a36e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h28f; din <= 32'hc6ef0ec4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h364; din <= 32'h96fb45a9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h010; din <= 32'h7049434f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h136; din <= 32'h43015f29;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h232; din <= 32'ha61e9045;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h197; din <= 32'hb2416b80;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h30a; din <= 32'h98108511;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08f; din <= 32'he83543f8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h121; din <= 32'h77716dbe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31c; din <= 32'hab38846d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h148; din <= 32'he21f0046;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23d; din <= 32'h1f94649b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e3; din <= 32'h7691dee2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d4; din <= 32'h2a1ee9df;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b2; din <= 32'h284b0de2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h25d; din <= 32'h7dda39aa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0fd; din <= 32'h102685d9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h398; din <= 32'h1e55d7e8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1cb; din <= 32'h972cb70e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b0; din <= 32'hb97cc2c5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3fe; din <= 32'hf46f92e4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h172; din <= 32'hf6453ac4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h03f; din <= 32'h0eda9024;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h398; din <= 32'hc2cae487;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h004; din <= 32'h6e4ab81e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h26e; din <= 32'he9fa261f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h29d; din <= 32'h568ccb01;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h057; din <= 32'h709c40ae;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37d; din <= 32'h4057f515;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a3; din <= 32'h93934c28;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h10b; din <= 32'h3805d83c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a0; din <= 32'h28fba0c5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ef; din <= 32'h56fec098;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h12e; din <= 32'hb3474b43;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h11b; din <= 32'h2abb061e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ae; din <= 32'hda6af91d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h190; din <= 32'hc4d209d1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a0; din <= 32'h4aef456e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37c; din <= 32'h2312ef1a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h069; din <= 32'h2ed405f6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3cb; din <= 32'hf01a2143;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h014; din <= 32'hc8c6555c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h300; din <= 32'ha58552fe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ca; din <= 32'h4cba39ae;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ec; din <= 32'h3d65e25d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b8; din <= 32'h6fe35927;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h17d; din <= 32'h8574ab9c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h136; din <= 32'h3c6f049f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h01a; din <= 32'h90dc2dbd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00f; din <= 32'h22ccbcf7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h10d; din <= 32'h69c2616b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ee; din <= 32'h7fc4683a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h203; din <= 32'h4169372a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2bd; din <= 32'h72b96d33;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h30a; din <= 32'h888a4ea9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h094; din <= 32'hd5356a57;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22d; din <= 32'h67c6ec8d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h35b; din <= 32'he5a16f20;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h390; din <= 32'h9aab446b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h192; din <= 32'h8287a37b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f2; din <= 32'hdb454610;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h06b; din <= 32'hdc8838ca;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c3; din <= 32'h22899408;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ae; din <= 32'h5eb6a999;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h396; din <= 32'h7344c334;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h21f; din <= 32'hd2a0ffb6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38b; din <= 32'hdcb10709;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h022; din <= 32'hcc3ce65f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h265; din <= 32'h683f2d5e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h09b; din <= 32'h00112435;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3fb; din <= 32'ha8e41a7c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h266; din <= 32'h854c8e0b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c9; din <= 32'h00e3974f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23b; din <= 32'h74c326ec;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0bb; din <= 32'h04f3bbed;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h25c; din <= 32'h05d0dc7d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h17e; din <= 32'hd3a67268;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1cb; din <= 32'h036f6e12;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h074; din <= 32'h27076e1a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h016; din <= 32'h2ecedf6d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h178; din <= 32'h29809773;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h21b; din <= 32'hf86e0e06;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c1; din <= 32'hf7c79a9a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h370; din <= 32'hcbc7d4ba;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e6; din <= 32'h1b8555d4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f0; din <= 32'h2f346fa2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h301; din <= 32'h186f17c3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h01a; din <= 32'h81b992f0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ef; din <= 32'h4f57c319;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3bf; din <= 32'ha5efccbb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h12d; din <= 32'hbec89bdf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h338; din <= 32'h9ab1cbc2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e6; din <= 32'hd5337799;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h07e; din <= 32'h61c9676a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h008; din <= 32'h3c5a332c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22e; din <= 32'h216657bf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f8; din <= 32'hbceab7a3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h168; din <= 32'h5a21f438;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c6; din <= 32'h30269070;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3db; din <= 32'hefcf664c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h248; din <= 32'hef39a5cc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f3; din <= 32'h6beefd0f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h20b; din <= 32'hdcdff49e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h063; din <= 32'h8dc3d16e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h303; din <= 32'h80fd3ede;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2cb; din <= 32'hbcb2e21a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h01b; din <= 32'h638585a9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h105; din <= 32'h043ffe2e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a9; din <= 32'hd4003647;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ec; din <= 32'hb24d0247;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h256; din <= 32'hac034b5a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h347; din <= 32'hc7ed9a43;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f5; din <= 32'h06457a19;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h020; din <= 32'hd18b24be;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h096; din <= 32'h041651e1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h11e; din <= 32'ha3ddc7a3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d9; din <= 32'h6d79ab91;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h398; din <= 32'hcb230c31;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1fa; din <= 32'h9525cc4b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d8; din <= 32'hdfdff08a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16a; din <= 32'h7f7d9a9a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ce; din <= 32'hf95b46a8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h398; din <= 32'h52ab10e2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h14f; din <= 32'h8f5f438b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h024; din <= 32'h12d2f99b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c4; din <= 32'he84a0b47;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2be; din <= 32'h075aa510;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b7; din <= 32'hc9891860;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h062; din <= 32'hf45e5ba3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c6; din <= 32'h513801df;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h30e; din <= 32'h4e203003;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h06c; din <= 32'h4eb61c68;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0be; din <= 32'hdac4099e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h021; din <= 32'h5b98ec72;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f4; din <= 32'h9681cc2d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h054; din <= 32'h4d3bb40b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f9; din <= 32'h8be31f8e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h002; din <= 32'h9ac2f15c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h190; din <= 32'h550b22cf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h222; din <= 32'h3c0ca15c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h064; din <= 32'h8a05bc7d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h32a; din <= 32'hc1882dba;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h068; din <= 32'hddaec768;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ce; din <= 32'h1527d925;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h13f; din <= 32'h6a236994;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h231; din <= 32'hfbe94a9a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h097; din <= 32'hd35ca39a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h227; din <= 32'h1eabed50;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h257; din <= 32'ha70524b1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h004; din <= 32'h5a88c87c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c1; din <= 32'h5441a34d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h27d; din <= 32'h8bd5174a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22f; din <= 32'h5710f167;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h13e; din <= 32'h74a66c7d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f2; din <= 32'h7c9c1514;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ba; din <= 32'hd318c8e8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c6; din <= 32'h9c10f096;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h284; din <= 32'hc3b22ea4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h350; din <= 32'h84a90557;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h220; din <= 32'h74525d69;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31c; din <= 32'h1f2fc523;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2a0; din <= 32'h277ddb7b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a0; din <= 32'h84e81735;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h034; din <= 32'h253dbc7e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2a8; din <= 32'h6d7a2813;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b3; din <= 32'h10d2edb9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ed; din <= 32'h18978809;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c0; din <= 32'h76d6bad6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h33b; din <= 32'h039b5c0f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h010; din <= 32'hecb0c960;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f7; din <= 32'h86ce63e1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d9; din <= 32'h07df22e5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d9; din <= 32'h7ab45dd8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h227; din <= 32'h6dce773b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h362; din <= 32'hd869136b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16e; din <= 32'ha562cb31;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c3; din <= 32'h06626513;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h356; din <= 32'hdce85a08;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h231; din <= 32'h3dac927f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e2; din <= 32'h75c80d91;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b8; din <= 32'h63cbcbaf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f9; din <= 32'h11c6aeb0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h09d; din <= 32'h6ae005b0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h352; din <= 32'hac67b187;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2aa; din <= 32'he5f11be5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e2; din <= 32'he6c0849e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h006; din <= 32'h07722846;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c7; din <= 32'ha9f753ca;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h034; din <= 32'h7c1ca9e1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0de; din <= 32'h03794b1c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h216; din <= 32'hb452f30d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h09b; din <= 32'ha74ad370;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f7; din <= 32'hedd4412a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18c; din <= 32'heb9347b5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h146; din <= 32'h224ec025;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h24a; din <= 32'hb90f6a53;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d4; din <= 32'h6e1d2c9d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d6; din <= 32'h8595ed1c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0cd; din <= 32'hb388e58f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h06e; din <= 32'h48c067f5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0fe; din <= 32'hb4e47fee;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a6; din <= 32'hcb4b0641;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h32b; din <= 32'hd43ae4b5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3af; din <= 32'he9a54d62;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h279; din <= 32'hc8b1fbf7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f2; din <= 32'h07b51fc9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h34a; din <= 32'h5cc24276;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h380; din <= 32'h70c5bce1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h353; din <= 32'h2c5d58c6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16b; din <= 32'h2b6c0293;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h028; din <= 32'hd289d15b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c5; din <= 32'hfd90435b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h30c; din <= 32'hcb20ff48;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a7; din <= 32'hd3e23302;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h17b; din <= 32'h4eb80889;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h234; din <= 32'h670b1c9d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h335; din <= 32'h7ed6252c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3bc; din <= 32'hd09b90d3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22f; din <= 32'h1c549b99;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b1; din <= 32'h92affa50;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c6; din <= 32'h74d6f74e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c4; din <= 32'hf7cb688b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b7; din <= 32'h918ecc39;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0bb; din <= 32'h59daee81;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h19c; din <= 32'h4ea3d581;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h19b; din <= 32'h2092ad67;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h01f; din <= 32'hdf3a45e5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a5; din <= 32'hf0f7f93a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h108; din <= 32'h28b7bf60;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ad; din <= 32'had084c8b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h073; din <= 32'h8ca6a013;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h061; din <= 32'h9c3953e7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d2; din <= 32'hbcc8fc88;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h338; din <= 32'h758efa46;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h20d; din <= 32'h364604db;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1bb; din <= 32'hb1328303;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h279; din <= 32'h030f9b41;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h32c; din <= 32'h5c748c0c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h199; din <= 32'h5de6e9fb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h088; din <= 32'h38be9c07;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h05a; din <= 32'h2fa02bb4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h089; din <= 32'hf5a54008;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h26f; din <= 32'he6aff25b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h309; din <= 32'h92015813;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h15e; din <= 32'hac95d379;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2cd; din <= 32'haed253b7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h20c; din <= 32'h5210c8ec;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18c; din <= 32'he5106006;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h197; din <= 32'h78cbb7e9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f4; din <= 32'heab748e0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h106; din <= 32'h013f8474;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h122; din <= 32'h7333a892;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d4; din <= 32'hcd129742;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16d; din <= 32'hbf13a884;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b8; din <= 32'he4b7b0ba;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h177; din <= 32'h04787c56;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h15c; din <= 32'h8e9f50b7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h34b; din <= 32'hd80f73ee;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h101; din <= 32'hf5753cc2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h062; din <= 32'h1b0bc678;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h042; din <= 32'hbb424e2b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h264; din <= 32'h3aa4372e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h074; din <= 32'hd72faebf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c3; din <= 32'h5d7d3855;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h119; din <= 32'ha0464d3e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00f; din <= 32'hfa7651d5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h224; din <= 32'h1f2c57a7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h343; din <= 32'hd23c83cf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h025; din <= 32'h3289dc51;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22d; din <= 32'ha1ec5eaf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f8; din <= 32'hb1c3ae7e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h214; din <= 32'h74948209;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h347; din <= 32'hececba0d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h125; din <= 32'h298eafa5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h05e; din <= 32'h696a928f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h368; din <= 32'h55a32397;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c0; din <= 32'hc1773d48;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f4; din <= 32'h832728c1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h13c; din <= 32'h2e59b6d8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ab; din <= 32'hd85cb9ae;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37e; din <= 32'h08dada69;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d3; din <= 32'he9c5599f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f5; din <= 32'h58c713e1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h262; din <= 32'hb842b354;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f8; din <= 32'h329703eb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h303; din <= 32'hd545bd0a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h284; din <= 32'h00a73ad5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f0; din <= 32'h1356e500;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f5; din <= 32'h9180cd99;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ab; din <= 32'heb6c11de;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h181; din <= 32'h2e9184bb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h368; din <= 32'hea45733f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h10e; din <= 32'h05a585bf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h052; din <= 32'h9436cb40;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h063; din <= 32'hae63e1a9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2cc; din <= 32'he566234d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h164; din <= 32'h15327b71;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h060; din <= 32'h38b9fce3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b2; din <= 32'hbedae9b2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e4; din <= 32'hee38965f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h074; din <= 32'hede615af;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ac; din <= 32'h0f604db8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2aa; din <= 32'h7e9ae6df;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h183; din <= 32'hd64e9fb3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b4; din <= 32'ha967896d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d1; din <= 32'h054a35bf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h130; din <= 32'hab5b8056;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h093; din <= 32'h5414f615;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d1; din <= 32'h33dd12dd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h175; din <= 32'h642f5a6c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h031; din <= 32'he8838bc0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h160; din <= 32'h6e741014;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a8; din <= 32'he94d299a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3dc; din <= 32'h4e90a475;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f9; din <= 32'h707ebba4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h029; din <= 32'h813be716;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3da; din <= 32'h4a611a2b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ad; din <= 32'h72b53f46;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h190; din <= 32'hb5751d6f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h079; din <= 32'h20a7ae45;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h241; din <= 32'hf634ecd4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ba; din <= 32'h39aefda9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h15e; din <= 32'h1e9ad03d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1fd; din <= 32'hc327343a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h191; din <= 32'hdaa3828b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b6; din <= 32'hd82d22b7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b5; din <= 32'h19c6dd8c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h28c; din <= 32'hc838403e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h216; din <= 32'h95a53430;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e5; din <= 32'hbaebe413;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h066; din <= 32'h9dba0923;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h03a; din <= 32'h969eb667;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31e; din <= 32'hbfe6e825;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0dc; din <= 32'h8760c752;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h329; din <= 32'h5ef4fa8e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h07a; din <= 32'h0c9510ed;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h149; din <= 32'h076e7536;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h025; din <= 32'h7a1d25ec;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d6; din <= 32'h42990661;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e7; din <= 32'h617a4d32;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h05b; din <= 32'h7943bf6b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2dc; din <= 32'h89d2be59;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31f; din <= 32'h2c967100;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a2; din <= 32'hb487ba2f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h153; din <= 32'h6e7b2a17;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38a; din <= 32'h63145bac;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1aa; din <= 32'h8dc077e8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b9; din <= 32'hbcc2164f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h251; din <= 32'ha7b26a87;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h174; din <= 32'h9e837615;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h032; din <= 32'hcb806db2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h19b; din <= 32'hb00061ce;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h17b; din <= 32'h3ff9d6b7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f8; din <= 32'h97cfafa1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22b; din <= 32'h8103a18e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h065; din <= 32'h165accaf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f2; din <= 32'hfdb67867;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e4; din <= 32'h412e4918;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h160; din <= 32'h078e289d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h165; din <= 32'h0559056b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b9; din <= 32'h5df7b0a6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h06a; din <= 32'hf48d9319;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h02b; din <= 32'h5026e52c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b7; din <= 32'hb241ddd0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h05e; din <= 32'h90acbcd2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h24a; din <= 32'he49483a9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a8; din <= 32'hcec4dde4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e6; din <= 32'h8ac7f211;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0fe; din <= 32'h439ad725;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h032; din <= 32'hc1a7ab81;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0af; din <= 32'h92c8c461;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3cd; din <= 32'h577cdaa0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h13d; din <= 32'hce5a3e59;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h025; din <= 32'h462db00f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h141; din <= 32'h28ed69d2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c6; din <= 32'h9eddae27;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3da; din <= 32'h44695257;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h013; din <= 32'h9b9a59d0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h215; din <= 32'h5a26da9f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h39e; din <= 32'h608e793a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h35e; din <= 32'hed037aaa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h20e; din <= 32'h13b3fa72;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h022; din <= 32'h37f033be;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ee; din <= 32'h5c55d30c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h192; din <= 32'hc37a0664;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a6; din <= 32'hd3dfd554;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h088; din <= 32'h1110396a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h296; din <= 32'h780b2dff;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h170; din <= 32'h4d883de7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h285; din <= 32'h557d4378;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h125; din <= 32'h7e4a75f6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h05c; din <= 32'h7ddc4274;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h02f; din <= 32'h0cfcc166;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h051; din <= 32'hdc8bfaaf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e6; din <= 32'h7dbe9b66;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h186; din <= 32'h46f8bb23;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ec; din <= 32'h6701567b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h29b; din <= 32'h7c4ed029;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h288; din <= 32'h86b7ff07;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h265; din <= 32'hec36df7f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h03a; din <= 32'h2f1fc535;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d4; din <= 32'hd378c891;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h13a; din <= 32'h5ef7ed16;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h073; din <= 32'h05616d2c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16a; din <= 32'hec0e01ff;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h125; din <= 32'heb6f7cf9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h003; din <= 32'h3e597b34;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h02b; din <= 32'hf4ced945;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h352; din <= 32'h028ddc3a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h197; din <= 32'h5549ccdd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ee; din <= 32'h54d08cff;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h12f; din <= 32'h348e3221;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c3; din <= 32'h22188188;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h12d; din <= 32'hec67aae5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f4; din <= 32'h7d2f6471;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h09b; din <= 32'h85b01651;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h024; din <= 32'hb35a0c85;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c9; din <= 32'h14d2d001;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h29d; din <= 32'hf3cfb48b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h34d; din <= 32'hdea2c3ff;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c6; din <= 32'h2dccbd0c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h332; din <= 32'hae583b60;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h110; din <= 32'hb2c10182;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h11e; din <= 32'hc4274337;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31a; din <= 32'h5179cbb8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b1; din <= 32'h5fa0e09e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h331; din <= 32'h2b121c79;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f5; din <= 32'hecf39c04;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ad; din <= 32'h758881bc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h228; din <= 32'h87e2e356;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h051; din <= 32'hd377030b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e5; din <= 32'h96a4c204;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d2; din <= 32'h51aee505;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c5; din <= 32'h71173c9d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h159; din <= 32'h2995928b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h030; din <= 32'h8c8bbb32;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31d; din <= 32'h30dfddd2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f7; din <= 32'he7d3077e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h124; din <= 32'h57888919;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h26f; din <= 32'hcc283f52;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h220; din <= 32'hb08656f1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ab; din <= 32'hfcea1007;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e2; din <= 32'h291b6884;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h013; din <= 32'hcd820473;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h11e; din <= 32'hb152407f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f4; din <= 32'h3ec0d07e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h342; din <= 32'h2a0d62fc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h152; din <= 32'hb89cdd2e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1df; din <= 32'hbbf94621;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h13a; din <= 32'hfe9f0a4e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e6; din <= 32'hbe615be4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h135; din <= 32'haec61891;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d2; din <= 32'hc260acda;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h34a; din <= 32'h6f9f6520;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h122; din <= 32'h8f2fba49;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h340; din <= 32'hc29471d7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37f; din <= 32'hed909107;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c3; din <= 32'hd9c3feb7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e3; din <= 32'h87f646b6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h016; din <= 32'h3cfdeafe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h27b; din <= 32'h589aeee4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h03e; din <= 32'h66d4f709;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a1; din <= 32'h91928457;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h32f; din <= 32'h78657504;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h390; din <= 32'he72df277;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1cf; din <= 32'h62eefe1f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ee; din <= 32'h01f78383;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h369; din <= 32'hbcac0dc8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3aa; din <= 32'h7f147473;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e9; din <= 32'ha0aeaf54;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h327; din <= 32'haf0e969f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h39f; din <= 32'h18dd8fd6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c3; din <= 32'hece70f5a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b4; din <= 32'h12e5061d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e4; din <= 32'he36e8757;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0db; din <= 32'h6b59e841;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h191; din <= 32'h7f4134db;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h102; din <= 32'h02fa04e8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2fd; din <= 32'hd2c1448b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1bd; din <= 32'h972d46af;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0cb; din <= 32'hc6f00bad;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h29d; din <= 32'h79b221e1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c4; din <= 32'haba3f8b6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0fe; din <= 32'h58d485bb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h240; din <= 32'hdaa1da74;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2dc; din <= 32'h77377687;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h224; din <= 32'h2537144e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b2; din <= 32'h35b51266;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h036; din <= 32'h7dbb491b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08f; din <= 32'hc31101f9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h159; din <= 32'hfe5d3235;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h125; din <= 32'hc3e5d8f8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b2; din <= 32'he42206e9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h186; din <= 32'hd90b6a14;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18d; din <= 32'h97b44f20;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ce; din <= 32'h859e5d0b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1cd; din <= 32'hfb67c0c4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h285; din <= 32'hae04fe57;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h132; din <= 32'h08b379b8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h35c; din <= 32'he4d6bf43;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h29d; din <= 32'h46db38bd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h040; din <= 32'hc6a8605d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c1; din <= 32'hf4f96654;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h087; din <= 32'h4debd5b7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b0; din <= 32'ha371bd8f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h255; din <= 32'h178201d2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h090; din <= 32'h876d5e4a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h247; din <= 32'hfc50d1b4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h13c; din <= 32'h8a91f41a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e7; din <= 32'haf6ce98a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f4; din <= 32'h6596e843;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h183; din <= 32'h01cefdb9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h21a; din <= 32'hc88f479c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e5; din <= 32'hf956fa21;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h33b; din <= 32'h65ecdf68;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h144; din <= 32'hdbb74eb7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c1; din <= 32'hf5648345;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h26f; din <= 32'hb0704715;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h047; din <= 32'hb8df8d8f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h046; din <= 32'h1c6efa8a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h25d; din <= 32'hc5df1eba;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0db; din <= 32'h5aa555de;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h336; din <= 32'h26fe6b32;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ac; din <= 32'hdea93abd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ce; din <= 32'hfc626eed;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d1; din <= 32'h99f17888;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h236; din <= 32'h74c2ff2e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37e; din <= 32'h2f62f972;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23e; din <= 32'hd4229241;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h176; din <= 32'hd64a651a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h353; din <= 32'h6e32eecc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h30e; din <= 32'h3df55cc4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d8; din <= 32'ha73ed0c6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e8; din <= 32'h9fc0198c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h398; din <= 32'h695e2def;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h303; din <= 32'hee877a01;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h17e; din <= 32'h63b6a8a1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h308; din <= 32'h1df87159;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f5; din <= 32'h1cb1683f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h276; din <= 32'h40e823fa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h30a; din <= 32'hf9fd2d62;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f8; din <= 32'h7d6f3968;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2a2; din <= 32'h09726fd2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37e; din <= 32'h2951c110;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h09b; din <= 32'h242e4c65;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h07d; din <= 32'h0e0cb601;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h21e; din <= 32'h73e66e7d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23b; din <= 32'h8d2315f5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h036; din <= 32'h71249e62;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e7; din <= 32'h210eeb2f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h131; din <= 32'h9ac5b9b6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h305; din <= 32'h65466386;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c7; din <= 32'h6d5eb7a5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a8; din <= 32'he231683a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d4; din <= 32'h140dd09e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h151; din <= 32'h76738709;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c6; din <= 32'h2cf5960a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h195; din <= 32'hbe403f7b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h189; din <= 32'h50bacce0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ef; din <= 32'h8ad282fe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d9; din <= 32'h39cb61b5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h289; din <= 32'hbe54ff00;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h100; din <= 32'h55dc04ea;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38f; din <= 32'h41475d05;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h20b; din <= 32'h891a781b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h15b; din <= 32'had1b1a35;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c3; din <= 32'hbbba2d4e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h204; din <= 32'hcbb6303b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e0; din <= 32'h6c9042d5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1dc; din <= 32'h0d9b71dd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1af; din <= 32'hc5a7d46c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h07b; din <= 32'h024de5d1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h086; din <= 32'hf45cb8a5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h304; din <= 32'h57253b25;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c5; din <= 32'h3def359f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h346; din <= 32'he6600ec0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h03a; din <= 32'he4655459;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ae; din <= 32'had636079;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h321; din <= 32'h7f4229cf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h32a; din <= 32'h7de322ac;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h02b; din <= 32'h4d7f1ec0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h050; din <= 32'he625abae;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08e; din <= 32'hd223c242;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h365; din <= 32'haa55c661;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h081; din <= 32'h73300d3e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h13b; din <= 32'h017bf1a7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h003; din <= 32'hadab46ec;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h09e; din <= 32'ha8ea94d6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h01b; din <= 32'hafab0131;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1eb; din <= 32'ha7c978a8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h370; din <= 32'hdd0a0696;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h015; din <= 32'h38e6b8e7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h216; din <= 32'heef4d8db;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h398; din <= 32'hf6279fac;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22e; din <= 32'hd2c33486;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h075; din <= 32'h393ef3ce;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b1; din <= 32'h79ec2fea;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h285; din <= 32'hb4b8281d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38e; din <= 32'hfdb0307b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h245; din <= 32'h2339594e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d7; din <= 32'hebba1873;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38e; din <= 32'h73eff0eb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h398; din <= 32'h7f638125;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0db; din <= 32'ha8ed1c06;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h326; din <= 32'h4bce0fa3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h103; din <= 32'h6a815f55;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h123; din <= 32'hb54acf26;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f9; din <= 32'h02f43054;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h280; din <= 32'h807b024c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c2; din <= 32'heb255876;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a4; din <= 32'hdfac93b5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h063; din <= 32'h32ef65dc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h131; din <= 32'h263ab781;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h210; din <= 32'hfa802e46;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b8; din <= 32'h7ef97a9b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h35e; din <= 32'h0730ae33;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h279; din <= 32'h1ca88af2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b0; din <= 32'hb2107507;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ea; din <= 32'hc6ae610d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b4; din <= 32'hbeb97d65;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h396; din <= 32'ha8c0f142;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b2; din <= 32'h5ffedba9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h36d; din <= 32'he0df0d82;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d0; din <= 32'h4a9e3b4c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d5; din <= 32'h8c71c29e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h106; din <= 32'he3f1d805;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d1; din <= 32'h3792b2cf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h19f; din <= 32'h7083fae5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16e; din <= 32'hc8cd1663;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h06a; din <= 32'h63eb66b9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d5; din <= 32'h0cf8cd51;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h357; din <= 32'h94733999;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f2; din <= 32'h0943ccea;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h321; din <= 32'hf1ad0a7e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h287; din <= 32'h8f272b08;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e0; din <= 32'h1f33dbae;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h337; din <= 32'hb73151a2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h255; din <= 32'h08e75b8b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22f; din <= 32'h2949684b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h279; din <= 32'h0b98b2b5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16d; din <= 32'h2874f9db;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h185; din <= 32'h682e08fb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h002; din <= 32'hac4e0b9e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h20a; din <= 32'h8ee28c40;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c2; din <= 32'hbccae8ad;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h048; din <= 32'h0b03ddc8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h135; din <= 32'h3a58125f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h19b; din <= 32'h430c6d81;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ef; din <= 32'hdef1c8fd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h36b; din <= 32'h7a516d0e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h10d; din <= 32'h8d4d88e0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h078; din <= 32'h0b364f94;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3fa; din <= 32'hdfd9e52c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2af; din <= 32'h32811267;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h379; din <= 32'hded09029;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1fd; din <= 32'h3a08452e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e2; din <= 32'hbd22fb13;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ee; din <= 32'h6575c8ab;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h13e; din <= 32'h8373ab10;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c8; din <= 32'hcc9a8907;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h318; din <= 32'h3ec9b6db;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h17e; din <= 32'hd501f135;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h10d; din <= 32'hdd68b8b1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h374; din <= 32'hb4fd02cb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h373; din <= 32'h57fcc8b3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h03d; din <= 32'h19a0e410;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0cc; din <= 32'hb338a54d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22a; din <= 32'h51bcab46;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b9; din <= 32'h97916cd1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h19c; din <= 32'h751fb28b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h203; din <= 32'hba332fb1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a6; din <= 32'h04608ed3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1dc; din <= 32'h8a5e68e7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h298; din <= 32'hfc3db7fa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h232; din <= 32'hcaee45f7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1de; din <= 32'hd3048179;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e0; din <= 32'h0cf7fdd5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h028; din <= 32'ha49e7716;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a7; din <= 32'h38649b9d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h14c; din <= 32'h2c80bba3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h171; din <= 32'h763790a5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1db; din <= 32'ha7a083fa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08b; din <= 32'h42faa88e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h347; din <= 32'h0fba2eb5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37e; din <= 32'h454e8360;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h25b; din <= 32'h954a58e9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c8; din <= 32'h598236d4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h089; din <= 32'h5b285a4e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h085; din <= 32'h8be80a7b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ef; din <= 32'hc5a51e85;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2cb; din <= 32'h974b29c0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h031; din <= 32'h93b45f22;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h081; din <= 32'hdd0a2f62;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2af; din <= 32'hbf6de63a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b9; din <= 32'h5fedc3de;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3db; din <= 32'h1de29d7a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e3; din <= 32'h74489252;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h30c; din <= 32'h8d1433c5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h182; din <= 32'h77bf8dc0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h044; din <= 32'hd68b9a51;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h380; din <= 32'h3037d9f2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f1; din <= 32'hf375498a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h262; din <= 32'ha817d4a8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h34a; din <= 32'ha962a302;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h311; din <= 32'h902fcb3a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c7; din <= 32'hb0e2e122;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h138; din <= 32'h6abc7b6e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h387; din <= 32'h6fbfdb9f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h14a; din <= 32'h2dd52a68;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h226; din <= 32'h08944558;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h30f; din <= 32'h56078150;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3af; din <= 32'hb239bf4f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h373; din <= 32'h0cbe1d63;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h138; din <= 32'h245ef888;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e3; din <= 32'h21c4382f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h077; din <= 32'hf4e829af;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2c7; din <= 32'h94cbd3ac;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22d; din <= 32'hf171bd32;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b5; din <= 32'he3d102ce;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h342; din <= 32'h0b1bc518;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f1; din <= 32'h41123bbb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h331; din <= 32'h0c9d146f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h04e; din <= 32'h71e6b58a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h185; din <= 32'had671e03;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h14b; din <= 32'h962f0a6a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h133; din <= 32'h044279b6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h379; din <= 32'h71ce9f89;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h235; din <= 32'he570d91a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h303; din <= 32'hf5dd0528;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h267; din <= 32'hc4e74286;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h25a; din <= 32'h1c78424c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h28d; din <= 32'h4e84674b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d1; din <= 32'hf6ecf4c1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d0; din <= 32'h7c5f15cd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h268; din <= 32'h7dfbc9ee;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h114; din <= 32'hf87b83f3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h280; din <= 32'h1253a283;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b6; din <= 32'hd2045758;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h153; din <= 32'hcc597153;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h208; din <= 32'h03660ebc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h330; din <= 32'h495cb63a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a4; din <= 32'h4691f4b1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h172; din <= 32'h81b0dd7f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f0; din <= 32'h907a8bf0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e3; din <= 32'h3abfec0b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ed; din <= 32'h1d2bd070;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b8; din <= 32'hd41bcdd1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h123; din <= 32'h03cca0b4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h33a; din <= 32'h9a97f30d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e6; din <= 32'h29ada1dc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h010; din <= 32'ha802bf5c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h34d; din <= 32'hf1ae66c7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ca; din <= 32'hceac49d5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c4; din <= 32'hcf6ab42d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h07f; din <= 32'h90727072;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h15a; din <= 32'h142b57a3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c2; din <= 32'hfb728343;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f2; din <= 32'heab7db96;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h185; din <= 32'hff416a36;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h10a; din <= 32'h39cecd56;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c4; din <= 32'h19f1bd04;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h276; din <= 32'h7fabd987;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3db; din <= 32'hd2f93e28;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h331; din <= 32'hdca18175;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h251; din <= 32'h888ff762;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h252; din <= 32'h5324c512;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h288; din <= 32'h0ad104d3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38a; din <= 32'hfa1816df;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h227; din <= 32'h4f2e7663;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23f; din <= 32'h06a49d2c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h038; din <= 32'hedb1f78a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d8; din <= 32'h46a7da5d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3fb; din <= 32'hd505998d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h180; din <= 32'hd0658924;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h379; din <= 32'h71130b5b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31b; din <= 32'h47c97b10;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h15c; din <= 32'h9bd00135;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37d; din <= 32'hf547798b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h054; din <= 32'he77dd1f5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h033; din <= 32'h17421646;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h233; din <= 32'h7c75ccbe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f2; din <= 32'h5512de86;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h076; din <= 32'hdde6a02b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h244; din <= 32'h64036466;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h338; din <= 32'h92f1773d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1fc; din <= 32'h4aa1a35e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b4; din <= 32'hd10afcc9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h25a; din <= 32'h9e92cc3f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h14c; din <= 32'h57e7c13f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h380; din <= 32'hd0a6db8a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c8; din <= 32'h6229fccb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f3; din <= 32'h798e0226;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h392; din <= 32'h54284ad7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h03e; din <= 32'hce786bf2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d6; din <= 32'h67e65135;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f6; din <= 32'h0c4cc681;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38b; din <= 32'h93f2925d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h318; din <= 32'h667c4f06;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d5; din <= 32'h91fa19ff;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d7; din <= 32'h50306075;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ad; din <= 32'hd8a775f3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h197; din <= 32'hb5c1c822;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h27e; din <= 32'ha5acaf94;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0bb; din <= 32'hd6fa2fcc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ca; din <= 32'ha52fdfc7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b4; din <= 32'hc0174ffe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h291; din <= 32'h06b37088;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h223; din <= 32'h538999f2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h352; din <= 32'h9adc7cd5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h039; din <= 32'h4e55e823;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h10a; din <= 32'hef802ad7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h178; din <= 32'hbbb979fa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b7; din <= 32'ha9aa3c64;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h157; din <= 32'h79dcfd08;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h318; din <= 32'h86ca738e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18e; din <= 32'h45e0ffe2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18b; din <= 32'hee1dee30;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h048; din <= 32'h19668afa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c0; din <= 32'h9bf8398d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d3; din <= 32'h4349a736;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h026; din <= 32'h26a10f85;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ad; din <= 32'h229e95bc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h256; din <= 32'h24c98b46;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16b; din <= 32'h6e3acbb3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h02c; din <= 32'h1e86147b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1bb; din <= 32'h349dbb46;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0e1; din <= 32'h86c95c9a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h289; din <= 32'h468ca22a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e1; din <= 32'hb606c33e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h395; din <= 32'hf0e89a2b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b2; din <= 32'hd84ccee8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h18a; din <= 32'h6c5efafd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f1; din <= 32'h528692b2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h013; din <= 32'h2521dd9c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h301; din <= 32'h1c199b3c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h211; din <= 32'h176c13c9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h12c; din <= 32'hc72c4364;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f8; din <= 32'h1dba2879;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b7; din <= 32'h8d41c3f6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h25f; din <= 32'hbbaa2b6e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a8; din <= 32'hf1d14ba1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f6; din <= 32'h4b13ba62;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h391; din <= 32'h488f81ec;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h34a; din <= 32'haedc68e2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h212; din <= 32'h2868bca6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h068; din <= 32'hfdd5cdb3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h098; din <= 32'hd0a88a76;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h186; din <= 32'h53b13a53;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b8; din <= 32'hae3b0212;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e6; din <= 32'h11d1be4a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f4; din <= 32'h3946c2fe;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h361; din <= 32'h7e1b51d8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h04d; din <= 32'h04e40c3d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h032; din <= 32'hce689197;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h373; din <= 32'h03846105;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h024; din <= 32'h257275d3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h35b; din <= 32'hf626449e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f1; din <= 32'h0ac68aaf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h03b; din <= 32'h5f1af0bd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h244; din <= 32'hdb578251;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h170; din <= 32'he8280dd1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0f4; din <= 32'h0294f659;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h07f; din <= 32'h98cac2e3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h239; din <= 32'h25524f48;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2df; din <= 32'h095a2e33;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h261; din <= 32'he621a0e9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d2; din <= 32'h1f419dcd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h28e; din <= 32'ha5cb5334;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e8; din <= 32'h1e823cbd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h162; din <= 32'h5661ff0f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22e; din <= 32'hcb29add1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1bd; din <= 32'hd3127b2f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f9; din <= 32'h34be2230;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2a5; din <= 32'h56dc2573;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h28b; din <= 32'hf92759c3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h266; din <= 32'h73ad522f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h072; din <= 32'hd9002dbd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h128; din <= 32'h25c7d640;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h341; din <= 32'he15e11a6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e4; din <= 32'h6b339af5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h087; din <= 32'hfd03cc03;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h05a; din <= 32'hbe8b2f5a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b0; din <= 32'h5eb0b5aa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h333; din <= 32'hf2d981c2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1bc; din <= 32'h6aae1902;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h002; din <= 32'h5eea5842;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h14e; din <= 32'h83d0eb90;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h07f; din <= 32'h9d7d45e7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ed; din <= 32'h95c3bc07;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b7; din <= 32'h2f0329d7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h06f; din <= 32'h9b0cfb2d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h215; din <= 32'hff43eb12;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c5; din <= 32'h775ee8b6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h045; din <= 32'hc1f2ff3c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b7; din <= 32'h74ee386b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h210; din <= 32'hd7ad697d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f9; din <= 32'h6a1e294a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h04e; din <= 32'h9848b616;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00f; din <= 32'h53dc1a30;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0de; din <= 32'h8ad319c4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37c; din <= 32'hfffd96be;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2a2; din <= 32'hafb05a84;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h21b; din <= 32'h26d4234f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31d; din <= 32'h25edb7a8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h219; din <= 32'h7bf87cb0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b6; din <= 32'h7500cd34;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h32a; din <= 32'h29337cc8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h11e; din <= 32'h7fc9c6ee;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h021; din <= 32'h7a3b6f3c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h120; din <= 32'hd1feddcb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h17b; din <= 32'h80f65570;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ae; din <= 32'h7339d19d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h241; din <= 32'h7b42a2b8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h194; din <= 32'hf3aa8e5b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h21e; din <= 32'h9a2c6864;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ae; din <= 32'h53b4fb83;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h13b; din <= 32'h4424f655;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h224; din <= 32'h647e73a5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b1; din <= 32'hde1eb12a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h227; din <= 32'h02944b17;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h130; din <= 32'h40b4e918;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h39b; din <= 32'h503d9ab7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h292; din <= 32'h6b9f1b5c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h32c; din <= 32'h494e0350;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h000; din <= 32'hb06f7d52;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h132; din <= 32'hd532829a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h297; din <= 32'h46adeff0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1a1; din <= 32'hcd53762d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ee; din <= 32'h9afed595;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h352; din <= 32'hd2b8f9f1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h13b; din <= 32'h29ca234f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2a9; din <= 32'h024a2777;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h238; din <= 32'h5c2e6d8e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a7; din <= 32'h921b6e79;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c7; din <= 32'hbc049ab9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h133; din <= 32'hc082ec61;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h278; din <= 32'hc3903ae6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h33b; din <= 32'h92a64bd6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h233; din <= 32'h26b6362f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h207; din <= 32'hd35ce640;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h048; din <= 32'hceeeae44;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c4; din <= 32'h71fa9986;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h308; din <= 32'ha4e98ade;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c2; din <= 32'hd5d29802;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h38a; din <= 32'haac0c56d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h11e; din <= 32'h0446a029;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h267; din <= 32'h5021d202;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0a6; din <= 32'hb0d3e5e3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0fc; din <= 32'h182f11f0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h01e; din <= 32'h15d22d32;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h36f; din <= 32'ha87095a5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h17c; din <= 32'h16d9d7ca;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b9; din <= 32'h8501bfbf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h381; din <= 32'h4ef6717b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f7; din <= 32'h335e6709;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0de; din <= 32'h5648cfa3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c2; din <= 32'hea1a0a80;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h15a; din <= 32'hd5b6a8c1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h35c; din <= 32'hf331bfbf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h395; din <= 32'hc3ae248a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d0; din <= 32'h30d403d0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1af; din <= 32'hb4fbd1dc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f6; din <= 32'h278c1c9f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h204; din <= 32'h5d1c46de;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h17b; din <= 32'hd38f592a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3b6; din <= 32'h76a6ee92;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16a; din <= 32'h65a8b943;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h363; din <= 32'h1bcb80da;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ee; din <= 32'h268ea449;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h380; din <= 32'h0de0fd9a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a5; din <= 32'hadf84edf;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h355; din <= 32'h6fdb06e4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d6; din <= 32'ha604825e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h33c; din <= 32'h4759ff22;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d7; din <= 32'h87b2aea5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h382; din <= 32'h00f4d630;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h291; din <= 32'h5e378bb8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h157; din <= 32'h66ad5c67;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c3; din <= 32'h63cd90da;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h324; din <= 32'hd24f77aa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h276; din <= 32'hd46e29c0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h313; din <= 32'h1b8147d5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h218; din <= 32'hd6e4059b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h320; din <= 32'hf927dcd5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ba; din <= 32'h38a1b16f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h045; din <= 32'hf1af31c8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h139; din <= 32'heaa4dd10;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h216; din <= 32'h560a6a66;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h332; din <= 32'h56644b1f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h141; din <= 32'h6c86dbb3;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23e; din <= 32'h87cb8c46;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3df; din <= 32'hc18ea6e1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h013; din <= 32'h8d16b057;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h393; din <= 32'h44c61ca2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1e1; din <= 32'hb44c37f6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h128; din <= 32'h4834b186;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h07e; din <= 32'h3eb27361;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d9; din <= 32'h837a0595;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h087; din <= 32'h0342ce34;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3d8; din <= 32'hb4293db6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ab; din <= 32'h4fb631b6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b6; din <= 32'hb83760ee;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d6; din <= 32'h6c3ca1e1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0bf; din <= 32'h3a14a624;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h065; din <= 32'he98cad7d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b1; din <= 32'h4f8be4f9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h127; din <= 32'heef3770c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h232; din <= 32'hb345bb00;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h193; din <= 32'hf704f3e4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h20f; din <= 32'h320bd0f6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h389; din <= 32'h1bb2b585;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ce; din <= 32'hf02e1867;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h116; din <= 32'h081306ea;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3aa; din <= 32'h868c242c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h33b; din <= 32'h01bdea60;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ff; din <= 32'hc64a02ff;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2d8; din <= 32'h836b5564;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1c6; din <= 32'head6f453;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h300; din <= 32'hcedfed04;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0c8; din <= 32'h3616a382;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h122; din <= 32'h636d4557;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h24d; din <= 32'hab4f1680;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b5; din <= 32'h7052d204;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h279; din <= 32'h7f411661;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h03e; din <= 32'h5d2fa9af;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h163; din <= 32'h2f89162b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h08f; din <= 32'h01605111;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h11b; din <= 32'hcf50681e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h24f; din <= 32'h88403ab8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1d3; din <= 32'h97a945d2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h19f; din <= 32'h2b7384a0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h26e; din <= 32'h95b13cbc;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22c; din <= 32'h7ce810aa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h235; din <= 32'h6ee41dfa;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h29a; din <= 32'hba79f510;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e8; din <= 32'h6695af01;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h14a; din <= 32'he8693b8f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e4; din <= 32'hcb818113;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h302; din <= 32'h2527ef95;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0aa; din <= 32'hbd89bc12;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h37b; din <= 32'h4258221b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h207; din <= 32'h89ad3fdd;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h050; din <= 32'he480e5e2;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h393; din <= 32'hee72768e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h287; din <= 32'h15c6a306;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2f2; din <= 32'h708467e4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h26b; din <= 32'ha1b3135e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1df; din <= 32'h5d863c19;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h154; din <= 32'hec64d91a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h21e; din <= 32'hc28095ac;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2ee; din <= 32'h9037e0c1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e9; din <= 32'h3f9ceeb5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h145; din <= 32'hb0a96673;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h27f; din <= 32'h7fb7182f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b6; din <= 32'h4dfe6b9d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h100; din <= 32'h251b2080;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h395; din <= 32'h713c64b4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h19d; din <= 32'hd5b94360;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h114; din <= 32'ha3ffd811;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h351; din <= 32'h2cf2939d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h090; din <= 32'h16279f1f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h329; din <= 32'h6f93878a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h22d; din <= 32'h7b3ba30d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h087; din <= 32'hed49cd4c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h184; din <= 32'h402c2aa7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f4; din <= 32'hc1ac3072;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h357; din <= 32'ha5d7f5f7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h00f; din <= 32'h984e4e1d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h374; din <= 32'h0ca5b8bb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e7; din <= 32'h208009a8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h237; din <= 32'hed0229b9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h195; din <= 32'h699020df;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e0; din <= 32'hcc436f2b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h14d; din <= 32'he91ed0d0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h298; din <= 32'he2829769;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h102; din <= 32'h6654048f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ff; din <= 32'h1d646100;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2b7; din <= 32'h46c9ab3f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h200; din <= 32'h2f79c051;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h16c; din <= 32'h5d394ef6;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h287; din <= 32'hdc786c0a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h095; din <= 32'h02955684;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0d5; din <= 32'h21215317;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h334; din <= 32'h988e9d9f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h241; din <= 32'h3fb03cad;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h21e; din <= 32'ha43796f1;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h108; din <= 32'h7268df91;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3eb; din <= 32'h4f6735d9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h13c; din <= 32'he85f458f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h33d; din <= 32'h35119895;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h36f; din <= 32'h17a03d53;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1ff; din <= 32'hc8ad01bb;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h23c; din <= 32'h78518d21;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h06a; din <= 32'h1b389e30;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h34c; din <= 32'h03230296;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h210; din <= 32'hf9505c38;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h214; din <= 32'h759c75d7;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1f2; din <= 32'h12c5fad8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h080; din <= 32'heef27a26;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h30c; din <= 32'ha25888c4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h29a; din <= 32'h07927808;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b8; din <= 32'h97d60f44;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h167; din <= 32'h9147b812;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h14b; din <= 32'ha9f5d670;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0ad; din <= 32'h77bf9d41;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h31e; din <= 32'h65256d26;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h062; din <= 32'h4cbd0a0f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3a3; din <= 32'h7511c352;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h0b0; din <= 32'hcc369a06;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h24f; din <= 32'h8a68fe5e;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h227; din <= 32'h9b076eb4;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h372; din <= 32'h5e3744e5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3fb; din <= 32'hc1bd269c;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1b2; din <= 32'h8fbf6c46;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h174; din <= 32'h4758283f;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h315; din <= 32'h71c1be0a;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h193; din <= 32'hc57b4f90;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e8; din <= 32'h98576f7b;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e6; din <= 32'h868214c5;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h184; din <= 32'hd4b9083d;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3e1; din <= 32'h5b0d08df;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3ac; din <= 32'h53891114;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3c4; din <= 32'h57737db0;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h319; din <= 32'h9d1848e8;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h1dc; din <= 32'h51820b38;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h118; din <= 32'h819b7cde;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h2e7; din <= 32'h6eaaeae9;
        @(posedge clk); op <= `NO_INSTR; addr <= 10'h3f6; din <= 32'he02e3cf4;

        // Finish
        @(posedge clk); op <= `NO_INSTR; addr <= 10'hxxx; din <= 32'hxxxxxxxx;
        repeat (5) @(posedge clk);
        $finish();
    end

    always #1 clk = ~clk;
endmodule
